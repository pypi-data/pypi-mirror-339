netcdf data {
dimensions:
	time = UNLIMITED ; // (15 currently)
variables:
	float time(time) ;
		time:unit = "s" ;
		time:label = "time" ;
	int STEP(time) ;
		STEP:label = "Palier" ;
	float PR1(time) ;
		PR1:unit = "bar" ;
		PR1:label = "PR1S" ;
	float PR15(time) ;
		PR15:unit = "bar" ;
		PR15:label = "PR15S" ;
	float PR30(time) ;
		PR30:unit = "bar" ;
		PR30:label = "PR30S" ;
	float PR60(time) ;
		PR60:unit = "bar" ;
		PR60:label = "PR60S" ;
	float PG1(time) ;
		PG1:unit = "bar" ;
		PG1:label = "PG1S" ;
	float PG15(time) ;
		PG15:unit = "bar" ;
		PG15:label = "PG15S" ;
	float PG30(time) ;
		PG30:unit = "bar" ;
		PG30:label = "PG30S" ;
	float PG60(time) ;
		PG60:unit = "bar" ;
		PG60:label = "PG60S" ;
	float V1(time) ;
		V1:unit = "cm3" ;
		V1:label = "V1S" ;
	float V15(time) ;
		V15:unit = "cm3" ;
		V15:label = "V15S" ;
	float V30(time) ;
		V30:unit = "cm3" ;
		V30:label = "V30S" ;
	float V60(time) ;
		V60:unit = "cm3" ;
		V60:label = "V60S" ;
		V60:scale_max = 500.f ;
	float CREEP(time) ;
		CREEP:unit = "cm3" ;
		CREEP:label = "fluage" ;
	float DELT60(time) ;
		DELT60:unit = "cm3" ;
		DELT60:label = "delt60" ;
data:

 time = 80, 141, 204, 269, 332, 398, 462, 525, 588, 652, 715, 778, 842, 906, 
    973 ;

 STEP = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 PR1 = 0.05, 0.88, 1.83, 3.02, 3.82, 8.73, 13.15, 17.69, 22.39, 26.94, 31.48, 
    36.02, 40.73, 45.42, 49.99 ;

 PR15 = 0.06, 0.81, 1.83, 2.95, 3.82, 8.5, 13.06, 17.68, 22.25, 26.81, 31.42, 
    36.07, 40.68, 45.32, 49.76 ;

 PR30 = 0.04, 0.82, 1.81, 2.95, 3.83, 8.48, 13.1, 17.69, 22.28, 26.82, 31.45, 
    36.06, 40.74, 45.36, 49.78 ;

 PR60 = 0.06, 0.82, 1.83, 2.93, 3.84, 8.48, 13.08, 17.72, 22.29, 26.84, 
    31.46, 36.11, 40.7, 45.31, 49.76 ;

 PG1 = 0.1, 0.11, 0.78, 1.82, 2.83, 7.37, 12.02, 16.69, 21.17, 25.89, 30.39, 
    35.01, 39.64, 44.37, 48.74 ;

 PG15 = 0.11, 0.08, 0.79, 1.81, 2.81, 7.39, 12.04, 16.61, 21.14, 25.77, 30.4, 
    35.01, 39.62, 44.29, 48.65 ;

 PG30 = 0.12, 0.11, 0.79, 1.81, 2.78, 7.41, 12, 16.61, 21.15, 25.78, 30.41, 
    35.02, 39.66, 44.31, 48.65 ;

 PG60 = 0.11, 0.09, 0.76, 1.8, 2.78, 7.37, 12.03, 16.65, 21.17, 25.8, 30.41, 
    35.04, 39.64, 44.28, 48.65 ;

 V1 = 31, 56, 168, 236, 240, 248, 250, 251, 253, 255, 255, 257, 257, 258, 259 ;

 V15 = 43, 98, 222, 237, 240, 247, 250, 251, 253, 254, 255, 257, 257, 258, 259 ;

 V30 = 46, 124, 229, 237, 240, 247, 249, 252, 253, 254, 255, 256, 258, 258, 
    258 ;

 V60 = 49, 152, 230, 238, 240, 247, 250, 252, 253, 254, 255, 257, 258, 258, 
    259 ;

 CREEP = 3, 28, 1, 1, 0, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1 ;

 DELT60 = 49, 103, 78, 8, 2, 7, 3, 2, 1, 1, 1, 2, 1, 0, 1 ;
}
