netcdf data {
dimensions:
	time = UNLIMITED ; // (42 currently)
variables:
	float time(time) ;
		time:unit = "s" ;
		time:label = "Temps" ;
	float DEPTH(time) ;
		DEPTH:unit = "m" ;
		DEPTH:label = "Prof." ;
	float AS(time) ;
		AS:unit = "m/h" ;
		AS:label = "VA" ;
		AS:scale_max = 800.f ;
	int EVP(time) ;
		EVP:label = "evt-part" ;
	int EVR(time) ;
		EVR:label = "evt-new-rod" ;
	float TP(time) ;
		TP:unit = "bar" ;
		TP:label = "PO" ;
		TP:scale_max = 200.f ;
	float IP(time) ;
		IP:unit = "bar" ;
		IP:label = "PI" ;
		IP:scale_max = 20.f ;
	float TQ(time) ;
		TQ:unit = "bar" ;
		TQ:label = "CR" ;
		TQ:scale_max = 200.f ;
	float SP(time) ;
		SP:unit = "bar" ;
		SP:label = "PF" ;
		SP:scale_max = 0.f ;
data:

 time = 0, 11.8, 12.6, 12.8, 13.8, 14, 14.2, 15.2, 15.4, 16, 16.2, 16.4, 
    16.8, 17.2, 17.4, 17.6, 17.8, 18.6, 19, 19.6, 20.2, 20.6, 21, 21.6, 22.2, 
    22.6, 23.2, 23.6, 24.2, 24.6, 25.2, 25.6, 26, 26.2, 26.4, 26.8, 27, 27.2, 
    27.4, 27.8, 48, 330.4 ;

 DEPTH = 0, 0.03, 0.04, 0.08, 0.09, 0.11, 0.12, 0.14, 0.16, 0.18, 0.2, 0.22, 
    0.23, 0.24, 0.27, 0.3, 0.32, 0.34, 0.36, 0.37, 0.38, 0.39, 0.4, 0.41, 
    0.42, 0.44, 0.45, 0.46, 0.47, 0.48, 0.5, 0.52, 0.53, 0.54, 0.55, 0.59, 
    0.6, 0.63, 0.65, 0.66, 0.68, 0.7 ;

 AS = 0.6613566, 8.576679, 45.18072, 686.747, 39.75904, 445.7831, 192.7711, 
    65.06024, 343.3735, 90.36144, 439.759, 391.5663, 93.3735, 99.39759, 
    463.8554, 524.0964, 421.6867, 91.86747, 147.5904, 60.24096, 60.24096, 
    93.3735, 93.3735, 68.27309, 80.32128, 117.4699, 76.30522, 90.36144, 
    60.24096, 111.4458, 86.34538, 180.7229, 99.39759, 216.8675, 277.1084, 
    280.1205, 331.3253, 457.8313, 409.6385, 105.4217, 3.459382, 6.024096 ;

 EVP = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EVR = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TP = 0, 62.35, 36.71, 73.34, 19.62, 66.01, 23.29, 70.89, 35.49, 9.86, 55.03, 
    79.44, 4.98, 14.74, 62.35, 78.22, 80.66, 46.48, 79.44, 79.44, 81.88, 
    81.88, 81.88, 81.88, 81.88, 79.44, 81.88, 81.88, 81.88, 81.88, 79.44, 
    81.88, 78.22, 78.22, 80.66, 80.66, 80.66, 80.66, 80.66, 70.89, 61.13, 0 ;

 IP = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TQ = 0, 78.22, 81.88, 81.88, 80.66, 80.66, 85.54, 80.66, 90.43, 90.43, 
    85.54, 89.21, 103.85, 95.31, 90.43, 97.75, 109.96, 111.18, 119.72, 
    124.61, 119.72, 113.62, 111.18, 105.07, 105.07, 109.96, 111.18, 111.18, 
    113.62, 113.62, 113.62, 125.83, 135.59, 138.03, 138.03, 130.71, 130.71, 
    128.27, 124.61, 150.24, 101.41, 0 ;

 SP = 661.72, 661.72, 661.72, 661.72, 661.72, 661.72, 661.72, 661.72, 661.72, 
    661.72, 661.72, 661.72, 661.72, 661.72, 661.72, 661.72, 661.72, 661.72, 
    661.72, 661.72, 661.72, 661.72, 661.72, 661.72, 661.72, 661.72, 661.72, 
    661.72, 661.72, 661.72, 661.72, 661.72, 661.72, 661.72, 661.72, 661.72, 
    661.72, 661.72, 661.72, 661.72, 661.72, 661.72 ;
}
