
module mod1;

    initial begin
        $display("mod1");
        $finish;
    end

endmodule
