netcdf data {
dimensions:
	time = UNLIMITED ; // (1203 currently)
variables:
	float time(time) ;
		time:unit = "s" ;
		time:label = "Temps" ;
	float DEPTH(time) ;
		DEPTH:unit = "m" ;
		DEPTH:label = "Prof." ;
	float AS(time) ;
		AS:unit = "m/h" ;
		AS:label = "VIA" ;
		AS:scale_max = 500.f ;
	int EVP(time) ;
		EVP:label = "evt-part" ;
	int EVR(time) ;
		EVR:label = "evt-new-rod" ;
	float TP(time) ;
		TP:unit = "bar" ;
		TP:label = "PO" ;
		TP:scale_max = 150.f ;
	float IP(time) ;
		IP:unit = "bar" ;
		IP:label = "PI" ;
		IP:scale_max = 50.f ;
	float TQ(time) ;
		TQ:unit = "bar" ;
		TQ:label = "CR" ;
		TQ:scale_max = 200.f ;
	float HP(time) ;
		HP:unit = "bar" ;
		HP:label = "PR" ;
		HP:scale_max = 0.f ;
data:

 time = 0, 2.8, 4, 5.4, 8, 11.4, 15.4, 19.4, 23, 26.8, 29.6, 31.6, 32.8, 
    34.6, 36.4, 38.2, 40.2, 42, 44, 45.8, 49.2, 53.4, 56.6, 59.8, 63, 65.8, 
    68.2, 70.4, 73.2, 75.6, 78.4, 81.4, 83.4, 85.4, 87.8, 90.4, 92.6, 95, 
    96.8, 99, 101.6, 104, 106.4, 108.8, 111.4, 115.2, 120.4, 125.2, 128.8, 
    133.2, 136, 139.2, 142.8, 146, 149, 152.8, 157.4, 162.2, 167.2, 172.6, 
    177, 181, 185.4, 189.8, 194.4, 199.4, 205, 210.2, 214.8, 218.4, 221, 
    222.6, 223.8, 226.6, 229.6, 233, 236.2, 239.6, 242.8, 246.4, 250, 253.8, 
    257.6, 261, 265.4, 269.6, 273.8, 277.8, 280.8, 283.6, 286.8, 290.2, 293, 
    296, 299, 302, 305.4, 308.6, 312.4, 316.2, 319.8, 323.4, 326.8, 329.6, 
    332, 333.8, 335.4, 337.2, 338.8, 340.6, 342.8, 344.8, 346.4, 348.6, 
    350.8, 353.8, 357.6, 361.4, 365.2, 368.2, 371.8, 376, 380.4, 384.2, 
    387.2, 390.4, 393.4, 395.2, 396.8, 399.2, 401.2, 404.4, 407.8, 412.2, 
    416.6, 420.6, 424.8, 428.2, 430.2, 431.8, 433.2, 434.8, 436.8, 439.6, 
    441.6, 443.8, 447, 451.6, 457.6, 462.6, 466, 468.6, 470.8, 473.2, 475.6, 
    478.8, 482.6, 486.6, 491.2, 494.8, 497.6, 499.6, 501, 502.4, 503.4, 
    504.4, 506, 509.4, 513.4, 516.599, 520.2, 522.8, 525.8, 528.6, 531, 
    533.6, 535.2, 537.2, 645.6, 647, 648.8, 650.4, 653.6, 655, 657, 658.6, 
    660.2, 662, 664.6, 667.8, 671.8, 674.6, 676.8, 679.8, 682.4, 684.4, 686, 
    687.6, 689, 690.4, 691.6, 692.8, 694, 695.4, 696.8, 700, 704, 708.8, 
    713.2, 717.6, 722, 724.6, 726.8, 729, 730.8, 732.2, 733.2, 734.2, 735, 
    736, 737, 738, 739, 740.2, 741.2, 742.2, 743.4, 744.6, 746, 747.8, 750, 
    752, 753.8, 755.6, 758.8, 763, 766.8, 769.6, 771.8, 773.6, 775.4, 778, 
    780.4, 782.4, 784.6, 786.8, 788.8, 790.6, 793.2, 796.4, 800.8, 804.6, 
    807, 808.6, 810.2, 811.6, 812.8, 814.4, 815.8, 817.4, 818.8, 820.2, 
    821.6, 823.2, 825, 827.2, 829.4, 832, 834.6, 837.2, 840, 843.6, 846.6, 
    849.4, 852.6, 855.4, 858, 861, 863.6, 865.6, 868, 871.4, 873.2, 875.6, 
    878.4, 881, 884.2, 886.4, 889.2, 892.2, 895, 898, 900.4, 903.4, 907, 910, 
    913.8, 917.2, 920.6, 924, 927, 931.2, 934.4, 938.4, 941.4, 944.4, 947.4, 
    950.4, 953.4, 956, 958.6, 961.4, 964, 967, 969.6, 972.4, 975, 977.4, 
    979.8, 982.2, 984.8, 987, 989.2, 991.8, 994, 996.6, 999, 1002, 1005.8, 
    1009, 1012.4, 1015.6, 1018.4, 1021.6, 1024.4, 1026.8, 1029.199, 1031.8, 
    1035, 1038.199, 1041.199, 1044, 1047, 1050.2, 1053, 1056.4, 1059, 1062, 
    1064.8, 1067.4, 1070.2, 1073, 1076, 1219, 1221.4, 1224, 1226.4, 1229, 
    1231.2, 1233.6, 1236, 1237.8, 1240, 1242, 1244.4, 1246.4, 1248, 1249.6, 
    1251, 1252.2, 1253.2, 1254.6, 1256.8, 1259, 1261.2, 1263.6, 1265.6, 
    1267.8, 1270.8, 1275.8, 1287.6, 1291.4, 1294.6, 1297.2, 1300.6, 1304.2, 
    1308.6, 1311.6, 1315.2, 1318.4, 1322.8, 1327.2, 1330, 1332.6, 1335.4, 
    1338, 1340.6, 1343, 1345.6, 1347.6, 1350.2, 1354.8, 1358.2, 1361.2, 
    1363.6, 1367.2, 1371.8, 1376.2, 1379.6, 1383.2, 1387.4, 1391.8, 1396.4, 
    1400.6, 1405, 1409.2, 1413.8, 1417.4, 1419.8, 1421.4, 1422.8, 1424, 
    1424.8, 1425.6, 1426.2, 1426.8, 1427.4, 1428, 1428.4, 1428.8, 1429.2, 
    1429.6, 1430.2, 1431.2, 1433.2, 1436.4, 1439.4, 1442.6, 1446.2, 1450, 
    1454, 1457.2, 1459.6, 1462.6, 1465.4, 1467.6, 1469.2, 1470.4, 1471.6, 
    1472.8, 1473.8, 1474.6, 1475.2, 1475.8, 1476.4, 1476.8, 1477.2, 1477.4, 
    1477.6, 1477.8, 1478, 1478.6, 1480.6, 1483.4, 1486.6, 1489.8, 1492.8, 
    1495.4, 1498, 1500.4, 1503, 1505.4, 1507.6, 1509.8, 1512.2, 1515, 1517.6, 
    1520.4, 1523.2, 1525.6, 1528.4, 1531.4, 1535, 1539.6, 1543.8, 1548.4, 
    1552.2, 1556.2, 1559.6, 1562.6, 1565.6, 1568, 1570, 1572.2, 1574.4, 
    1577.2, 1579.6, 1582.4, 1585.2, 1588.2, 1591.6, 1594.2, 1597.4, 1600.6, 
    1604.2, 1607.8, 1611, 1614.2, 1617.6, 1620.6, 1624.6, 1628, 1632, 1636, 
    1639.6, 1642.6, 1645.6, 1648.8, 1652, 1655.4, 1658.6, 1661.8, 1664.8, 
    1853.4, 1855.8, 1859, 1862, 1865.2, 1868.2, 1870.4, 1872.8, 1875.6, 
    1877.8, 1880.8, 1883.8, 1887.6, 1891.2, 1894.6, 1897.4, 1900.4, 1903.6, 
    1907, 1909.8, 1912.4, 1915.4, 1918.6, 1921.8, 1925.2, 1928.8, 1932.4, 
    1935.8, 1939, 1942, 1945.6, 1948.4, 1950.6, 1953.2, 1955.6, 1958.4, 1962, 
    1965.8, 1971, 1976.2, 1981, 1986, 1990.8, 1995.2, 1999.8, 2004.2, 2007.4, 
    2010.8, 2015, 2019, 2022.2, 2025, 2027.6, 2031.2, 2035.4, 2038.8, 2041.6, 
    2043.8, 2045.8, 2047.4, 2048.8, 2050.399, 2052.2, 2054.8, 2057, 2059, 
    2060.8, 2062.399, 2064.2, 2066.2, 2068.2, 2070.2, 2072.2, 2073.8, 2076, 
    2078.6, 2080.6, 2083, 2085.2, 2087.8, 2090.399, 2092.399, 2094.399, 
    2096.8, 2099.4, 2102.8, 2106.2, 2109.6, 2113.4, 2117, 2120.4, 2123.4, 
    2126.6, 2130.2, 2134.6, 2139.6, 2144.6, 2150.2, 2713.6, 2718.6, 2722.8, 
    2727, 2730.2, 2733.4, 2736.8, 2739.6, 2742.4, 2745, 2747.6, 2749.8, 2752, 
    2756, 2758.6, 2761.8, 2766.2, 2769.2, 2772.8, 2776.6, 2780.6, 2783.2, 
    2786.4, 2789.2, 2793.2, 2797.8, 2802.4, 2806.6, 2810.8, 2814.8, 2819, 
    2822.6, 2826.6, 2830.6, 2834.4, 2838.2, 2841.6, 2844.6, 2846.8, 2848.6, 
    2850.2, 2851.6, 2853.6, 2856.6, 2859.6, 2863.2, 2866.4, 2870.4, 2874.4, 
    2878, 2881.6, 2884, 2887.6, 2891.4, 2895.2, 2898.4, 2901.6, 2904.8, 
    2907.6, 2909.8, 2911.4, 2913.4, 2916.2, 2919, 2922.2, 2925.6, 2929, 
    2932.8, 2936.8, 2940.4, 2944, 2947.8, 2951.6, 2955.2, 2959, 2962.4, 2965, 
    2968.2, 2971.4, 2974.6, 2977.6, 2981, 2985, 2989, 2993.2, 2997.4, 3001.4, 
    3058.4, 3062.8, 3067, 3070.2, 3073, 3075.4, 3077, 3079.2, 3082, 3085, 
    3088.2, 3091.2, 3093.6, 3097, 3100.6, 3104.6, 3107, 3110, 3112.6, 3115.2, 
    3117.6, 3120.2, 3122.8, 3125.4, 3128.4, 3132.2, 3136, 3140, 3144.2, 
    3148.2, 3151.4, 3154.8, 3158.6, 3162, 3165.8, 3169.8, 3173.6, 3178.2, 
    3182.2, 3186.6, 3190.6, 3195, 3198.8, 3201, 3203.8, 3206.4, 3209.8, 
    3213.6, 3217.8, 3222.2, 3226.4, 3230.8, 3235.4, 3239.8, 3244.2, 3247.6, 
    3250.6, 3253.4, 3256.2, 3258.2, 3260.4, 3262, 3263.4, 3265.4, 3268.2, 
    3270.6, 3273, 3275.8, 3278.8, 3281.4, 3283.8, 3286.4, 3289.6, 3293, 
    3296.8, 3300.4, 3304.2, 3307.8, 3311.4, 3315.2, 3319, 3322.6, 3326.8, 
    3330.6, 3334.4, 3338, 3341.4, 3344.8, 3348.6, 3352.4, 3356.4, 3359.6, 
    3363, 3366.4, 3369.8, 3373.6, 3378, 3382, 3386, 3390, 3394.2, 3398.4, 
    3402.2, 3406.4, 3410.4, 3414.2, 3418, 3421.6, 3424.8, 3427.6, 3430, 
    3432.2, 3435, 3438.2, 3441.4, 3443.8, 3446.2, 3449.2, 3452.6, 3455, 
    3457.4, 3459.6, 3461.6, 3463.8, 3465.8, 3468, 3471, 3474.6, 3477.8, 
    3481.4, 3485, 3488.6, 3493, 3496.8, 3500.6, 3504.2, 3507.6, 3511.2, 
    3515.2, 3519.2, 3522.8, 3526.2, 3529.6, 3533.4, 3536.8, 3540.4, 3543.6, 
    3546.8, 3549.4, 3553.4, 3558, 3562.8, 3567.8, 3572, 3577, 3581, 3585.6, 
    3591, 3595.8, 3601.2, 3606.2, 3611.2, 3616.4, 3621, 3626, 3630.6, 3635.8, 
    3640.4, 3644.8, 3649.8, 3654.2, 3658.4, 3783.2, 3789, 3794.8, 3800.4, 
    3806, 3810.4, 3815.8, 3821, 3826.6, 3830.4, 3833.4, 3836.2, 3840.4, 
    3844.6, 3849.6, 3854.6, 3860, 3865.2, 3870.4, 3876, 3881.4, 3886.8, 3892, 
    3896.4, 3899, 3901.4, 3904, 3907.6, 3911.8, 3915.8, 3918.6, 3920.8, 
    3922.8, 3924.6, 3926.6, 3929.4, 3932.6, 3936, 3940, 3944.6, 3949, 3953.6, 
    3956.8, 3959.4, 3961.8, 3966.8, 3972.4, 3978.4, 3983.4, 3987.8, 3990.4, 
    3992, 3993.6, 3996.2, 4000, 4005.4, 4011, 4016.4, 4021.8, 4026.4, 4030.4, 
    4032.4, 4033.8, 4035.4, 4037.4, 4040.2, 4042.8, 4045.2, 4047.6, 4049.4, 
    4050.6, 4052.2, 4053.8, 4058, 4063.6, 4069.6, 4075, 4080.6, 4085.6, 
    4090.2, 4094.2, 4098, 4100, 4102, 4105.6, 4110.4, 4114.799, 4119.2, 
    4123.6, 4127.799, 4132.2, 4134.4, 4135.799, 4138, 4141.2, 4145, 4149.4, 
    4153.6, 4157.4, 4161.4, 4165.6, 4170, 4174.799, 4180.4, 4186.2, 4192, 
    4198, 4203.4, 4208.4, 4212, 4215, 4217.8, 4221, 4224.4, 4226.8, 4229.8, 
    4233, 4236.8, 4241.2, 4245.8, 4250, 4254.6, 4260, 4265.4, 4270.6, 4276, 
    4280.6, 4283.8, 4286.8, 4289.6, 4292.6, 4296.6, 4300.8, 4305.2, 4309.2, 
    4312.4, 4315.2, 4317.8, 4321.6, 4325.2, 4329.8, 4335.2, 4341, 4347.4, 
    4353.4, 4360, 4365.8, 4370.6, 4375, 4377.2, 4380.2, 4385.4, 4390.4, 4393, 
    4395, 4399, 4404, 4408.8, 4413.2, 4415.8, 4417.6, 4420.8, 4424.2, 4428.8, 
    4434, 4439.2, 4444.4, 4449.2, 4454.4, 4459, 4462.6, 4464.8, 4504, 4682.4, 
    4685.8, 4689, 4692.2, 4696, 4700.8, 4705, 4708.6, 4713.4, 4718.2, 4722.6, 
    4726, 4729.4, 4732.4, 4736.8, 4741.6, 4746.4, 4750.2, 4754.2, 4759.6, 
    4764.8, 4768.6, 4771.8, 4776.4, 4781, 4785.6, 4789.2, 4792, 4796.2, 
    4799.8, 4803, 4806, 4808.4, 4810.8, 4814.6, 4819.2, 4824, 4828, 4830.2, 
    4831.8, 4834.6, 4838.4, 4842.8, 4847.2, 4851.4, 4856, 4860, 4863.4, 
    4866.6, 4868.8, 4870.4, 4872.2, 4874.6, 4878.2, 4881.6, 4884.6, 4888, 
    4891.8, 4896, 4900.4, 4904.6, 4909, 4913.6, 4918.2, 4922.6, 4925.8, 
    4928.4, 4931, 4933, 4934.6, 4936.8, 4939.4, 4943.8, 4948.6, 4954.2, 
    4960.2, 4965, 4969.6, 4974, 4977.8, 4980.8, 4983.2, 4985, 4986.6, 4989, 
    4991.6, 4994.4, 4997, 4999.6, 5002.4, 5005.2, 5008.2, 5012, 5016.2, 
    5020.6, 5025.6, 5030, 5034.6, 5038.6, 5041.4, 5043.6, 5045, 5046, 5047.6, 
    5050, 5053.8, 5058.8, 5064, 5069.4, 5074.6, 5079, 5083, 5086.6, 5088.6, 
    5090.8, 5093.8, 5097.4, 5101.4, 5105.8, 5111, 5116.2, 5121.2, 5126.4, 
    5131.2, 5136.6, 5142, 5147.4, 5152, 5155.4, 5158.2, 5159.8, 5161.4, 
    5164.2, 5168.4, 5174.4, 5180.8, 5186.8, 5191.8, 5195.8, 5198.6, 5201.2, 
    5203, 5205.2, 5207.2, 5209, 5211.2, 5214, 5219.4, 5224.4, 5233.8 ;

 DEPTH = 7.71, 7.72, 7.73, 7.74, 7.75, 7.76, 7.77, 7.78, 7.79, 7.8, 7.81, 
    7.82, 7.83, 7.85, 7.86, 7.87, 7.88, 7.89, 7.9, 7.91, 7.92, 7.93, 7.94, 
    7.95, 7.96, 7.97, 7.98, 7.99, 8, 8.01, 8.02, 8.03, 8.04, 8.05, 8.06, 
    8.07, 8.08, 8.09, 8.1, 8.11, 8.12, 8.13, 8.14, 8.15, 8.16, 8.17, 8.18, 
    8.19, 8.2, 8.21, 8.22, 8.23, 8.24, 8.25, 8.26, 8.27, 8.28, 8.29, 8.3, 
    8.31, 8.32, 8.33, 8.34, 8.35, 8.36, 8.37, 8.38, 8.39, 8.4, 8.41, 8.42, 
    8.43, 8.44, 8.45, 8.47, 8.48, 8.49, 8.5, 8.51, 8.52, 8.53, 8.54, 8.55, 
    8.56, 8.57, 8.58, 8.59, 8.6, 8.61, 8.62, 8.63, 8.64, 8.65, 8.66, 8.67, 
    8.68, 8.69, 8.7, 8.71, 8.72, 8.73, 8.74, 8.75, 8.76, 8.77, 8.78, 8.79, 
    8.8, 8.81, 8.82, 8.83, 8.84, 8.85, 8.86, 8.87, 8.88, 8.89, 8.9, 8.91, 
    8.92, 8.93, 8.94, 8.95, 8.96, 8.97, 8.98, 8.99, 9, 9.01, 9.02, 9.03, 
    9.04, 9.05, 9.06, 9.07, 9.08, 9.09, 9.1, 9.11, 9.12, 9.14, 9.15, 9.16, 
    9.17, 9.18, 9.19, 9.2, 9.21, 9.22, 9.23, 9.24, 9.25, 9.26, 9.27, 9.28, 
    9.29, 9.3, 9.31, 9.32, 9.33, 9.34, 9.35, 9.36, 9.37, 9.38, 9.39, 9.4, 
    9.41, 9.42, 9.43, 9.44, 9.45, 9.46, 9.47, 9.48, 9.49, 9.5, 9.51, 9.52, 
    9.53, 9.54, 9.55, 9.57, 9.58, 9.59, 9.6, 9.61, 9.62, 9.63, 9.64, 9.65, 
    9.66, 9.67, 9.68, 9.69, 9.7, 9.71, 9.72, 9.73, 9.74, 9.75, 9.76, 9.77, 
    9.78, 9.79, 9.8, 9.81, 9.82, 9.83, 9.84, 9.85, 9.86, 9.87, 9.88, 9.89, 
    9.9, 9.91, 9.93, 9.94, 9.95, 9.96, 9.97, 9.98, 9.99, 10, 10.01, 10.02, 
    10.03, 10.04, 10.05, 10.06, 10.07, 10.08, 10.09, 10.1, 10.11, 10.12, 
    10.13, 10.14, 10.15, 10.16, 10.17, 10.18, 10.19, 10.2, 10.22, 10.23, 
    10.24, 10.25, 10.26, 10.27, 10.28, 10.29, 10.3, 10.31, 10.32, 10.33, 
    10.34, 10.35, 10.36, 10.37, 10.38, 10.39, 10.4, 10.41, 10.42, 10.43, 
    10.44, 10.45, 10.46, 10.47, 10.48, 10.49, 10.5, 10.51, 10.52, 10.53, 
    10.54, 10.56, 10.57, 10.58, 10.59, 10.6, 10.61, 10.62, 10.63, 10.64, 
    10.65, 10.66, 10.67, 10.68, 10.69, 10.7, 10.71, 10.72, 10.73, 10.74, 
    10.75, 10.76, 10.77, 10.78, 10.79, 10.8, 10.81, 10.82, 10.83, 10.84, 
    10.85, 10.86, 10.87, 10.88, 10.89, 10.9, 10.91, 10.92, 10.93, 10.94, 
    10.95, 10.96, 10.97, 10.98, 10.99, 11, 11.01, 11.02, 11.03, 11.04, 11.05, 
    11.06, 11.07, 11.08, 11.09, 11.1, 11.11, 11.12, 11.13, 11.14, 11.15, 
    11.16, 11.17, 11.18, 11.19, 11.2, 11.21, 11.22, 11.23, 11.24, 11.25, 
    11.26, 11.27, 11.28, 11.3, 11.31, 11.32, 11.33, 11.34, 11.35, 11.36, 
    11.37, 11.38, 11.39, 11.4, 11.41, 11.42, 11.43, 11.44, 11.45, 11.46, 
    11.47, 11.48, 11.49, 11.5, 11.51, 11.52, 11.53, 11.54, 11.55, 11.56, 
    11.57, 11.58, 11.59, 11.6, 11.61, 11.63, 11.64, 11.65, 11.66, 11.67, 
    11.68, 11.69, 11.7, 11.71, 11.72, 11.73, 11.74, 11.75, 11.76, 11.77, 
    11.78, 11.79, 11.8, 11.81, 11.82, 11.83, 11.84, 11.85, 11.86, 11.87, 
    11.88, 11.89, 11.9, 11.91, 11.92, 11.93, 11.94, 11.95, 11.96, 11.97, 
    11.98, 11.99, 12, 12.01, 12.02, 12.03, 12.05, 12.06, 12.07, 12.08, 12.09, 
    12.1, 12.11, 12.12, 12.13, 12.14, 12.15, 12.16, 12.17, 12.18, 12.19, 
    12.2, 12.22, 12.23, 12.24, 12.25, 12.26, 12.27, 12.28, 12.29, 12.3, 
    12.31, 12.32, 12.33, 12.34, 12.36, 12.37, 12.39, 12.4, 12.41, 12.42, 
    12.43, 12.44, 12.45, 12.47, 12.48, 12.49, 12.5, 12.51, 12.52, 12.53, 
    12.54, 12.55, 12.56, 12.57, 12.58, 12.59, 12.6, 12.61, 12.62, 12.63, 
    12.64, 12.65, 12.66, 12.67, 12.68, 12.69, 12.7, 12.71, 12.72, 12.73, 
    12.74, 12.75, 12.76, 12.77, 12.78, 12.79, 12.8, 12.81, 12.82, 12.83, 
    12.84, 12.85, 12.86, 12.87, 12.88, 12.89, 12.9, 12.91, 12.92, 12.93, 
    12.94, 12.95, 12.97, 12.98, 12.99, 13, 13.01, 13.02, 13.03, 13.04, 13.05, 
    13.06, 13.07, 13.08, 13.09, 13.1, 13.11, 13.12, 13.13, 13.14, 13.15, 
    13.16, 13.17, 13.18, 13.19, 13.2, 13.21, 13.22, 13.23, 13.24, 13.25, 
    13.26, 13.27, 13.28, 13.29, 13.3, 13.31, 13.32, 13.33, 13.34, 13.35, 
    13.36, 13.37, 13.38, 13.39, 13.4, 13.41, 13.42, 13.43, 13.44, 13.45, 
    13.47, 13.48, 13.49, 13.5, 13.51, 13.52, 13.53, 13.54, 13.55, 13.56, 
    13.57, 13.58, 13.59, 13.6, 13.61, 13.62, 13.63, 13.64, 13.65, 13.66, 
    13.67, 13.68, 13.69, 13.7, 13.71, 13.72, 13.73, 13.74, 13.75, 13.76, 
    13.77, 13.78, 13.79, 13.8, 13.81, 13.82, 13.83, 13.84, 13.85, 13.86, 
    13.88, 13.89, 13.9, 13.91, 13.92, 13.93, 13.94, 13.95, 13.96, 13.97, 
    13.98, 13.99, 14, 14.01, 14.02, 14.03, 14.04, 14.05, 14.06, 14.07, 14.08, 
    14.09, 14.1, 14.11, 14.12, 14.13, 14.14, 14.15, 14.16, 14.17, 14.18, 
    14.19, 14.2, 14.21, 14.22, 14.23, 14.24, 14.25, 14.26, 14.27, 14.28, 
    14.29, 14.3, 14.31, 14.32, 14.33, 14.34, 14.35, 14.36, 14.37, 14.38, 
    14.39, 14.4, 14.41, 14.42, 14.43, 14.44, 14.45, 14.47, 14.48, 14.49, 
    14.5, 14.51, 14.52, 14.53, 14.54, 14.55, 14.56, 14.57, 14.58, 14.59, 
    14.6, 14.61, 14.62, 14.63, 14.64, 14.65, 14.66, 14.67, 14.68, 14.69, 
    14.7, 14.71, 14.72, 14.73, 14.74, 14.75, 14.76, 14.77, 14.78, 14.79, 
    14.8, 14.81, 14.82, 14.83, 14.84, 14.85, 14.86, 14.87, 14.88, 14.89, 
    14.9, 14.91, 14.92, 14.93, 14.94, 14.95, 14.96, 14.97, 14.98, 14.99, 15, 
    15.01, 15.02, 15.04, 15.05, 15.06, 15.07, 15.08, 15.09, 15.1, 15.11, 
    15.12, 15.13, 15.14, 15.15, 15.16, 15.17, 15.18, 15.19, 15.2, 15.21, 
    15.22, 15.23, 15.24, 15.25, 15.26, 15.27, 15.28, 15.29, 15.3, 15.31, 
    15.32, 15.33, 15.34, 15.35, 15.36, 15.37, 15.38, 15.39, 15.4, 15.41, 
    15.42, 15.43, 15.44, 15.45, 15.46, 15.47, 15.48, 15.49, 15.5, 15.51, 
    15.52, 15.53, 15.54, 15.55, 15.56, 15.57, 15.58, 15.59, 15.6, 15.61, 
    15.63, 15.64, 15.65, 15.66, 15.67, 15.68, 15.69, 15.7, 15.71, 15.72, 
    15.73, 15.74, 15.75, 15.76, 15.77, 15.78, 15.79, 15.8, 15.81, 15.82, 
    15.83, 15.84, 15.85, 15.86, 15.87, 15.88, 15.89, 15.9, 15.91, 15.92, 
    15.93, 15.94, 15.95, 15.96, 15.97, 15.98, 15.99, 16, 16.01, 16.02, 16.03, 
    16.04, 16.05, 16.06, 16.07, 16.08, 16.09, 16.1, 16.11, 16.12, 16.13, 
    16.14, 16.15, 16.16, 16.17, 16.18, 16.19, 16.2, 16.21, 16.22, 16.23, 
    16.24, 16.25, 16.26, 16.27, 16.28, 16.29, 16.3, 16.31, 16.32, 16.33, 
    16.34, 16.35, 16.36, 16.38, 16.39, 16.4, 16.41, 16.42, 16.43, 16.44, 
    16.45, 16.46, 16.47, 16.48, 16.49, 16.5, 16.51, 16.52, 16.53, 16.54, 
    16.55, 16.56, 16.57, 16.58, 16.59, 16.6, 16.61, 16.62, 16.63, 16.64, 
    16.65, 16.66, 16.67, 16.68, 16.69, 16.7, 16.71, 16.72, 16.73, 16.74, 
    16.75, 16.76, 16.77, 16.78, 16.79, 16.8, 16.81, 16.82, 16.83, 16.84, 
    16.85, 16.86, 16.87, 16.88, 16.89, 16.9, 16.91, 16.92, 16.93, 16.94, 
    16.95, 16.97, 16.98, 16.99, 17, 17.01, 17.02, 17.03, 17.04, 17.05, 17.06, 
    17.07, 17.08, 17.09, 17.1, 17.11, 17.12, 17.13, 17.14, 17.15, 17.16, 
    17.17, 17.18, 17.19, 17.2, 17.21, 17.22, 17.23, 17.24, 17.25, 17.26, 
    17.27, 17.28, 17.29, 17.3, 17.31, 17.32, 17.33, 17.34, 17.35, 17.36, 
    17.37, 17.38, 17.39, 17.4, 17.41, 17.42, 17.43, 17.44, 17.45, 17.46, 
    17.47, 17.48, 17.49, 17.5, 17.51, 17.52, 17.53, 17.54, 17.55, 17.56, 
    17.57, 17.58, 17.59, 17.6, 17.61, 17.63, 17.64, 17.65, 17.66, 17.67, 
    17.68, 17.69, 17.7, 17.71, 17.72, 17.73, 17.74, 17.75, 17.76, 17.77, 
    17.78, 17.79, 17.8, 17.81, 17.82, 17.83, 17.84, 17.85, 17.86, 17.87, 
    17.88, 17.89, 17.9, 17.91, 17.92, 17.93, 17.94, 17.95, 17.96, 17.97, 
    17.98, 17.99, 18, 18.01, 18.02, 18.03, 18.04, 18.05, 18.06, 18.07, 18.08, 
    18.09, 18.1, 18.11, 18.12, 18.13, 18.14, 18.15, 18.16, 18.17, 18.18, 
    18.19, 18.2, 18.21, 18.22, 18.23, 18.24, 18.25, 18.26, 18.27, 18.28, 
    18.3, 18.31, 18.32, 18.33, 18.34, 18.35, 18.36, 18.37, 18.38, 18.39, 
    18.4, 18.41, 18.42, 18.43, 18.44, 18.45, 18.46, 18.47, 18.48, 18.49, 
    18.5, 18.51, 18.52, 18.53, 18.54, 18.55, 18.56, 18.57, 18.58, 18.59, 
    18.6, 18.61, 18.62, 18.63, 18.64, 18.65, 18.66, 18.67, 18.68, 18.69, 
    18.7, 18.71, 18.72, 18.73, 18.74, 18.75, 18.76, 18.77, 18.78, 18.79, 
    18.8, 18.81, 18.82, 18.83, 18.84, 18.85, 18.86, 18.87, 18.88, 18.89, 
    18.9, 18.91, 18.92, 18.93, 18.94, 18.95, 18.96, 18.97, 18.98, 18.99, 19, 
    19.01, 19.02, 19.03, 19.05, 19.06, 19.07, 19.08, 19.09, 19.1, 19.11, 
    19.12, 19.13, 19.14, 19.15, 19.16, 19.17, 19.18, 19.19, 19.2, 19.21, 
    19.22, 19.23, 19.24, 19.25, 19.26, 19.27, 19.28, 19.29, 19.3, 19.31, 
    19.32, 19.33, 19.34, 19.35, 19.36, 19.37, 19.38, 19.39, 19.4, 19.41, 
    19.42, 19.43, 19.44, 19.45, 19.46, 19.47, 19.48, 19.49, 19.5, 19.51, 
    19.52, 19.53, 19.54, 19.55, 19.56, 19.57, 19.58, 19.59, 19.6, 19.61, 
    19.62, 19.63, 19.64, 19.65, 19.66, 19.67, 19.68, 19.69, 19.7, 19.72, 
    19.73, 19.74, 19.75, 19.76, 19.77, 19.78, 19.79, 19.8, 19.81, 19.82, 
    19.83, 19.84, 19.85, 19.86, 19.87, 19.88, 19.89, 19.9, 19.91, 19.92, 
    19.93, 19.94, 19.95, 19.96, 19.97, 19.98, 20 ;

 AS = 0, 15.23161, 33.78378, 26.06178, 14.03326, 10.73132, 9.121622, 
    9.121622, 10.13513, 9.601707, 13.03089, 18.24324, 30.40541, 22.52252, 
    20.27027, 20.27027, 18.24324, 20.27027, 18.24324, 20.27027, 10.73132, 
    8.687259, 11.40203, 11.40203, 11.40203, 13.03089, 15.2027, 16.58477, 
    13.03089, 15.2027, 13.03089, 12.16216, 18.24324, 18.24324, 15.2027, 
    14.03326, 16.58477, 15.2027, 20.27027, 16.58477, 14.03326, 15.2027, 
    15.2027, 15.2027, 14.03326, 9.601707, 7.016632, 7.601351, 10.13513, 
    8.292383, 13.03089, 11.40203, 10.13513, 11.40203, 12.16216, 9.601707, 
    7.931845, 7.601351, 7.297297, 6.756757, 8.292383, 9.121622, 8.292383, 
    8.292383, 7.931845, 7.297297, 6.515444, 7.016632, 7.931845, 10.13513, 
    14.03326, 25.33784, 30.40541, 13.03089, 12.16216, 10.73132, 11.40203, 
    10.73132, 11.40203, 10.13513, 10.13513, 9.601707, 9.601707, 10.73132, 
    8.292383, 8.687259, 8.687259, 9.121622, 12.16216, 13.03089, 11.40203, 
    10.73132, 13.03089, 12.16216, 12.16216, 12.16216, 10.73132, 11.40203, 
    9.601707, 9.601707, 10.13513, 10.13513, 10.73132, 13.03089, 15.2027, 
    20.27027, 22.80405, 20.27027, 22.80405, 20.27027, 16.58477, 18.24324, 
    22.80405, 16.58477, 16.58477, 12.16216, 9.601707, 9.601707, 9.601707, 
    12.16216, 10.13513, 8.687259, 8.292383, 9.601707, 12.16216, 11.40203, 
    12.16216, 20.27027, 22.80405, 15.2027, 18.24324, 11.40203, 10.73132, 
    8.292383, 8.292383, 9.121622, 8.687259, 10.73132, 18.24324, 22.80405, 
    31.85328, 22.80405, 18.24324, 13.03089, 18.24324, 16.58477, 11.40203, 
    7.931845, 6.081081, 7.297297, 10.73132, 14.03326, 16.58477, 15.2027, 
    15.2027, 11.40203, 9.601707, 9.121622, 7.931845, 10.13513, 13.03089, 
    18.24324, 26.06178, 28.95753, 40.54054, 36.48649, 22.80405, 10.73132, 
    9.121622, 11.40203, 10.13513, 14.03326, 12.16216, 13.03089, 15.2027, 
    14.03326, 22.80405, 18.24324, 0.3365912, 26.06178, 20.27027, 22.80405, 
    12.66892, 26.06178, 18.24324, 22.80405, 22.80405, 20.27027, 14.03326, 
    11.40203, 9.121622, 13.03089, 16.58477, 12.16216, 15.59252, 18.24324, 
    22.80405, 22.80405, 28.95753, 26.06178, 30.40541, 30.40541, 30.40541, 
    28.95753, 26.06178, 11.40203, 9.121622, 7.601351, 8.292383, 8.292383, 
    8.292383, 14.03326, 16.58477, 16.58477, 20.27027, 26.06178, 36.48649, 
    44.59459, 45.60811, 36.48649, 40.54054, 36.48649, 36.48649, 33.78378, 
    36.48649, 40.54054, 33.78378, 30.40541, 26.06178, 20.27027, 16.58477, 
    18.24324, 20.27027, 20.27027, 11.40203, 8.687259, 9.601707, 13.03089, 
    16.58477, 20.27027, 20.27027, 15.59252, 15.2027, 18.24324, 16.58477, 
    16.58477, 18.24324, 20.27027, 14.03326, 11.40203, 8.292383, 9.601707, 
    15.2027, 22.80405, 22.80405, 26.06178, 30.40541, 25.33784, 26.06178, 
    25.33784, 26.06178, 26.06178, 26.06178, 22.80405, 20.27027, 16.58477, 
    16.58477, 14.03326, 14.03326, 14.03326, 13.03089, 10.13513, 12.16216, 
    13.03089, 11.40203, 13.03089, 15.59252, 13.51351, 15.59252, 18.24324, 
    15.2027, 10.73132, 20.27027, 15.2027, 13.03089, 14.03326, 11.40203, 
    16.58477, 13.03089, 12.16216, 13.03089, 12.16216, 15.2027, 12.16216, 
    10.13513, 12.16216, 9.601707, 10.73132, 10.73132, 10.73132, 12.16216, 
    8.687259, 11.40203, 9.121622, 12.16216, 12.16216, 12.16216, 12.16216, 
    12.16216, 14.03326, 14.03326, 13.03089, 14.03326, 12.16216, 14.03326, 
    13.03089, 14.03326, 15.2027, 15.2027, 15.2027, 14.03326, 16.58477, 
    16.58477, 14.03326, 16.58477, 14.03326, 15.2027, 12.16216, 9.601707, 
    11.40203, 10.73132, 11.40203, 13.03089, 11.40203, 13.03089, 15.2027, 
    15.2027, 14.03326, 11.40203, 11.40203, 12.16216, 13.03089, 12.16216, 
    11.40203, 13.03089, 10.73132, 14.03326, 12.16216, 13.03089, 14.03326, 
    13.03089, 13.03089, 12.16216, 0.2551503, 15.2027, 14.03326, 15.2027, 
    14.03326, 16.58477, 15.2027, 15.2027, 20.27027, 18.42752, 18.24324, 
    15.2027, 20.27027, 22.80405, 22.80405, 28.95753, 33.78378, 40.54054, 
    26.06178, 16.58477, 16.58477, 16.58477, 15.2027, 18.24324, 16.58477, 
    12.16216, 7.297297, 3.092075, 9.601707, 11.40203, 14.03326, 10.73132, 
    10.13513, 8.292383, 12.16216, 10.13513, 11.40203, 8.292383, 8.292383, 
    13.03089, 14.03326, 13.03089, 14.03326, 14.03326, 15.2027, 14.03326, 
    18.24324, 14.03326, 7.931845, 10.73132, 12.16216, 15.2027, 10.13513, 
    7.931845, 8.292383, 10.73132, 10.13513, 8.687259, 8.292383, 7.931845, 
    8.687259, 8.292383, 8.687259, 7.931845, 10.13513, 15.2027, 22.80405, 
    28.95753, 33.78378, 50.67567, 50.67567, 60.81081, 67.56757, 74.32433, 
    81.08108, 91.21622, 91.21622, 91.21622, 91.21622, 67.56757, 36.48649, 
    18.24324, 11.40203, 12.16216, 11.40203, 10.13513, 9.601707, 9.121622, 
    11.40203, 15.2027, 12.16216, 13.03089, 16.58477, 25.33784, 33.78378, 
    33.78378, 33.78378, 36.48649, 50.67567, 67.56757, 74.32433, 94.5946, 
    131.7568, 152.027, 182.4324, 182.4324, 182.4324, 182.4324, 67.56757, 
    18.24324, 13.03089, 11.40203, 11.40203, 12.16216, 14.03326, 14.03326, 
    15.2027, 14.03326, 15.2027, 16.58477, 16.58477, 15.2027, 13.03089, 
    14.03326, 13.03089, 13.03089, 15.2027, 13.03089, 12.16216, 10.13513, 
    7.931845, 8.687259, 7.931845, 9.601707, 9.121622, 10.73132, 13.51351, 
    13.51351, 15.2027, 18.24324, 16.58477, 18.42752, 13.03089, 15.2027, 
    13.03089, 13.03089, 12.16216, 10.73132, 14.03326, 11.40203, 11.40203, 
    10.13513, 10.13513, 11.40203, 11.40203, 10.73132, 12.16216, 9.121622, 
    10.73132, 9.121622, 9.121622, 10.13513, 12.16216, 12.16216, 11.40203, 
    11.40203, 10.73132, 11.40203, 11.40203, 12.16216, 0.1934596, 15.2027, 
    11.40203, 12.16216, 11.40203, 12.16216, 16.58477, 15.2027, 14.47876, 
    16.58477, 12.16216, 12.16216, 9.601707, 10.13513, 10.73132, 13.03089, 
    12.16216, 11.40203, 11.92369, 13.03089, 14.03326, 12.16216, 11.40203, 
    11.40203, 10.73132, 10.13513, 10.13513, 10.73132, 11.40203, 12.16216, 
    10.13513, 14.47876, 16.58477, 14.03326, 15.2027, 13.03089, 10.13513, 
    9.601707, 7.016632, 7.016632, 7.601351, 7.297297, 7.601351, 8.292383, 
    7.931845, 8.292383, 11.40203, 10.73132, 8.687259, 9.121622, 11.40203, 
    13.03089, 14.03326, 10.13513, 8.687259, 10.73132, 14.47876, 16.58477, 
    20.27027, 22.80405, 26.06178, 22.80405, 20.27027, 14.03326, 16.58477, 
    18.24324, 20.27027, 22.80405, 22.52252, 18.24324, 18.24324, 20.27027, 
    18.24324, 22.80405, 16.58477, 14.03326, 18.24324, 15.2027, 16.58477, 
    14.03326, 14.03326, 18.24324, 18.24324, 15.2027, 14.03326, 10.73132, 
    10.73132, 10.73132, 9.601707, 10.13513, 10.73132, 12.16216, 11.40203, 
    10.13513, 8.292383, 7.297297, 7.297297, 6.515444, 11.35144, 7.297297, 
    8.687259, 8.687259, 11.40203, 11.40203, 10.73132, 13.03089, 13.03089, 
    14.03326, 14.03326, 16.58477, 16.58477, 9.121622, 14.03326, 11.40203, 
    8.292383, 12.16216, 10.13513, 9.601707, 9.121622, 14.03326, 11.40203, 
    13.03089, 9.121622, 7.931845, 7.931845, 8.687259, 8.687259, 9.121622, 
    8.687259, 10.13513, 9.121622, 9.121622, 9.601707, 9.601707, 10.73132, 
    12.16216, 16.58477, 20.27027, 22.80405, 26.06178, 18.24324, 12.16216, 
    12.16216, 10.13513, 11.40203, 9.121622, 9.121622, 10.13513, 10.13513, 
    15.2027, 10.13513, 9.601707, 9.601707, 11.40203, 11.40203, 11.40203, 
    13.03089, 16.58477, 22.80405, 18.24324, 13.03089, 13.03089, 11.40203, 
    10.73132, 10.73132, 9.601707, 9.121622, 10.13513, 10.13513, 9.601707, 
    10.66856, 11.26126, 9.601707, 10.73132, 14.03326, 11.40203, 11.40203, 
    11.40203, 12.16216, 10.73132, 9.121622, 9.121622, 8.687259, 8.687259, 
    9.121622, 0.6401138, 8.292383, 8.687259, 11.40203, 13.03089, 15.2027, 
    25.33784, 16.58477, 13.03089, 12.16216, 11.40203, 12.16216, 15.2027, 
    10.73132, 10.13513, 9.121622, 15.2027, 12.16216, 14.03326, 14.03326, 
    15.2027, 14.03326, 14.03326, 14.03326, 12.16216, 9.601707, 9.601707, 
    9.121622, 8.687259, 9.121622, 11.40203, 10.73132, 9.601707, 10.73132, 
    9.601707, 9.121622, 9.601707, 7.931845, 9.121622, 8.292383, 9.121622, 
    8.292383, 9.601707, 16.58477, 14.47876, 14.03326, 10.73132, 9.601707, 
    8.687259, 8.292383, 8.687259, 8.292383, 7.931845, 8.292383, 8.292383, 
    10.73132, 12.16216, 13.03089, 13.03089, 18.24324, 16.58477, 22.80405, 
    26.06178, 18.24324, 13.03089, 15.2027, 15.2027, 13.03089, 12.16216, 
    14.03326, 15.2027, 14.03326, 11.40203, 10.73132, 9.601707, 10.13513, 
    9.601707, 10.13513, 10.13513, 9.601707, 9.601707, 10.13513, 8.687259, 
    9.601707, 9.601707, 10.13513, 10.73132, 10.73132, 9.601707, 9.601707, 
    9.121622, 11.40203, 10.73132, 10.73132, 10.73132, 9.601707, 8.292383, 
    9.121622, 9.121622, 9.121622, 8.687259, 8.687259, 9.601707, 8.687259, 
    9.121622, 9.601707, 9.601707, 10.13513, 11.40203, 13.03089, 15.2027, 
    16.58477, 13.03089, 11.40203, 11.40203, 15.2027, 15.2027, 12.16216, 
    10.73132, 15.2027, 15.2027, 16.58477, 18.24324, 16.58477, 18.24324, 
    16.58477, 12.16216, 10.13513, 11.40203, 10.13513, 10.13513, 10.13513, 
    8.292383, 9.601707, 9.601707, 10.13513, 10.73132, 10.13513, 9.121622, 
    9.121622, 10.13513, 10.73132, 10.73132, 9.601707, 10.73132, 10.13513, 
    11.40203, 11.40203, 14.03326, 9.121622, 7.931845, 7.601351, 7.297297, 
    8.687259, 7.297297, 9.121622, 7.931845, 6.756757, 7.601351, 6.756757, 
    7.297297, 7.297297, 7.016632, 7.931845, 7.297297, 7.931845, 7.016632, 
    7.931845, 8.292383, 7.297297, 8.292383, 8.687259, 0.2923597, 6.290773, 
    6.290773, 7.239382, 6.515444, 8.292383, 6.756757, 7.016632, 6.515444, 
    9.601707, 12.16216, 13.03089, 8.687259, 8.687259, 7.297297, 7.297297, 
    6.756757, 7.016632, 7.016632, 6.515444, 6.756757, 6.756757, 7.796258, 
    8.292383, 14.03326, 15.2027, 14.03326, 10.13513, 8.687259, 9.121622, 
    13.03089, 16.58477, 18.24324, 20.27027, 18.24324, 13.03089, 11.40203, 
    10.73132, 9.121622, 7.931845, 8.292383, 7.931845, 11.40203, 14.03326, 
    15.2027, 7.297297, 6.515444, 6.081081, 7.297297, 8.292383, 14.03326, 
    25.33784, 22.80405, 14.03326, 9.601707, 6.756757, 6.515444, 6.756757, 
    6.756757, 7.931845, 9.121622, 18.24324, 26.06178, 22.80405, 18.24324, 
    13.03089, 14.03326, 15.2027, 15.2027, 20.27027, 30.40541, 22.80405, 
    22.80405, 8.687259, 6.515444, 6.081081, 6.756757, 6.515444, 7.297297, 
    7.931845, 9.121622, 9.601707, 18.24324, 18.24324, 10.13513, 7.601351, 
    8.292383, 8.292383, 8.292383, 8.687259, 8.292383, 18.42752, 26.06178, 
    16.58477, 11.40203, 9.601707, 8.292383, 8.687259, 9.601707, 9.121622, 
    8.687259, 8.292383, 7.601351, 6.515444, 6.290773, 6.290773, 6.081081, 
    6.756757, 7.297297, 10.13513, 12.16216, 13.03089, 11.40203, 10.73132, 
    15.2027, 12.16216, 11.40203, 9.601707, 8.292383, 7.931845, 8.687259, 
    7.931845, 6.756757, 6.756757, 7.016632, 6.756757, 7.931845, 11.40203, 
    12.16216, 13.03089, 12.16216, 9.121622, 8.687259, 8.292383, 9.121622, 
    11.40203, 13.03089, 14.03326, 9.601707, 10.13513, 7.931845, 6.756757, 
    6.290773, 5.701014, 6.081081, 5.528255, 6.290773, 7.601351, 8.292383, 
    16.58477, 12.16216, 7.016632, 7.297297, 14.03326, 18.24324, 9.121622, 
    7.297297, 7.601351, 8.292383, 14.03326, 20.27027, 11.40203, 10.73132, 
    7.931845, 7.016632, 7.016632, 7.016632, 7.601351, 7.016632, 7.931845, 
    10.13513, 16.58477, 0.9307777, 0.2045207, 10.73132, 11.40203, 11.40203, 
    9.601707, 7.601351, 8.687259, 10.13513, 7.601351, 7.601351, 8.292383, 
    10.73132, 10.73132, 12.16216, 8.292383, 7.601351, 7.601351, 9.601707, 
    9.121622, 6.756757, 7.016632, 9.601707, 11.40203, 7.931845, 7.931845, 
    7.931845, 10.13513, 13.03089, 8.687259, 10.13513, 11.40203, 12.16216, 
    15.2027, 15.2027, 9.601707, 7.931845, 7.601351, 9.121622, 16.58477, 
    22.80405, 13.03089, 9.601707, 8.292383, 8.292383, 8.687259, 7.931845, 
    9.121622, 10.73132, 11.40203, 16.58477, 22.80405, 20.27027, 15.2027, 
    10.13513, 10.73132, 12.16216, 10.73132, 9.601707, 8.687259, 8.292383, 
    8.687259, 8.292383, 7.931845, 7.931845, 8.292383, 11.40203, 14.03326, 
    14.03326, 18.24324, 22.80405, 16.58477, 14.03326, 8.292383, 7.601351, 
    6.515444, 6.081081, 7.601351, 7.931845, 8.292383, 9.601707, 12.16216, 
    15.2027, 20.27027, 22.80405, 15.2027, 14.03326, 13.03089, 14.03326, 
    14.03326, 14.47876, 13.03089, 12.16216, 9.601707, 8.687259, 8.292383, 
    7.297297, 8.292383, 7.931845, 9.121622, 13.03089, 16.58477, 26.06178, 
    36.48649, 22.80405, 15.2027, 9.601707, 7.297297, 7.016632, 6.756757, 
    7.016632, 8.292383, 9.121622, 10.13513, 18.24324, 16.58477, 12.16216, 
    10.13513, 9.121622, 8.292383, 7.016632, 7.016632, 7.297297, 7.016632, 
    7.601351, 6.756757, 6.756757, 6.756757, 7.931845, 10.73132, 13.03089, 
    22.80405, 22.80405, 13.03089, 8.687259, 6.081081, 5.701014, 6.081081, 
    7.297297, 9.121622, 13.03089, 14.03326, 20.27027, 16.58477, 18.24324, 
    20.27027, 16.58477, 13.03089, 6.756757, 7.297297, 7.297297 ;

 EVP = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0 ;

 EVR = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0 ;

 TP = 53.2, 51.67, 51.67, 51.98, 51.98, 52.59, 52.59, 52.59, 52.59, 52.59, 
    52.28, 51.98, 51.98, 51.98, 51.67, 52.28, 52.59, 51.67, 52.28, 51.98, 
    51.98, 52.59, 51.98, 52.28, 52.28, 51.98, 51.98, 51.98, 51.67, 51.67, 
    51.67, 51.98, 51.67, 51.67, 51.98, 51.98, 51.67, 51.67, 51.67, 51.67, 
    51.98, 51.98, 51.67, 51.67, 51.98, 52.28, 52.28, 51.98, 52.28, 52.28, 
    52.28, 52.28, 51.98, 51.98, 51.98, 51.98, 52.28, 52.59, 54.72, 55.34, 
    54.72, 54.42, 55.03, 55.03, 55.03, 54.72, 54.42, 54.72, 55.03, 54.72, 
    54.42, 54.11, 54.11, 53.81, 54.72, 54.11, 53.81, 54.11, 54.42, 54.42, 
    54.42, 53.5, 54.72, 55.03, 54.72, 54.72, 54.42, 53.81, 54.11, 53.81, 
    53.81, 53.5, 53.2, 54.11, 54.42, 54.42, 54.42, 54.42, 54.42, 54.42, 
    54.72, 54.72, 54.42, 53.81, 54.42, 54.11, 54.11, 54.42, 54.11, 53.81, 
    54.11, 53.81, 54.42, 54.42, 54.11, 54.42, 54.42, 54.42, 53.5, 53.5, 
    54.42, 53.2, 54.72, 54.42, 53.5, 54.42, 54.11, 53.5, 53.5, 53.81, 53.81, 
    54.11, 54.42, 54.42, 54.11, 54.42, 53.81, 53.81, 54.11, 53.81, 52.59, 
    54.11, 54.11, 53.5, 53.81, 53.81, 54.11, 54.11, 53.5, 54.72, 54.11, 
    54.42, 54.42, 54.42, 54.72, 54.11, 54.72, 53.81, 54.42, 54.72, 54.11, 
    53.81, 53.5, 53.2, 53.5, 53.2, 54.42, 54.11, 53.81, 53.81, 53.5, 54.42, 
    54.42, 54.11, 54.11, 54.42, 53.81, 53.5, 53.81, 53.81, 53.5, 54.11, 
    52.28, 53.5, 53.5, 53.81, 54.11, 53.2, 54.42, 54.11, 53.81, 54.42, 54.42, 
    54.11, 53.5, 53.5, 53.5, 53.81, 53.2, 51.67, 51.37, 51.37, 51.37, 51.67, 
    51.37, 51.98, 51.98, 51.67, 51.67, 51.98, 51.98, 51.98, 52.28, 52.59, 
    52.89, 52.28, 51.98, 51.98, 52.28, 52.28, 51.67, 52.59, 52.59, 52.28, 
    51.98, 51.98, 52.28, 51.98, 52.28, 52.59, 52.59, 52.28, 52.59, 52.28, 
    52.59, 53.2, 52.89, 52.28, 52.28, 51.98, 52.59, 52.28, 51.98, 52.89, 
    52.28, 52.59, 52.28, 52.28, 52.59, 52.28, 52.59, 52.59, 52.28, 51.98, 
    52.28, 52.28, 52.59, 51.98, 51.98, 52.28, 51.67, 51.98, 52.28, 52.28, 
    52.28, 52.59, 52.59, 52.28, 52.59, 51.98, 52.28, 52.59, 52.28, 54.11, 
    55.34, 55.34, 55.64, 55.03, 55.34, 53.81, 55.64, 55.34, 55.34, 55.03, 
    55.03, 55.34, 53.2, 53.2, 53.2, 53.2, 52.89, 52.89, 52.89, 52.89, 52.28, 
    53.2, 53.2, 52.89, 53.2, 53.2, 52.89, 53.2, 53.2, 53.2, 52.89, 53.2, 
    52.89, 52.89, 52.28, 52.89, 52.89, 53.2, 53.2, 52.89, 52.89, 52.89, 
    52.59, 52.59, 52.89, 53.2, 52.59, 52.59, 52.28, 52.59, 52.59, 52.89, 
    52.28, 52.59, 52.89, 52.59, 52.89, 53.2, 53.2, 53.2, 52.59, 52.89, 52.59, 
    51.98, 53.2, 52.89, 52.89, 52.59, 52.89, 51.98, 52.89, 52.89, 52.89, 
    53.2, 53.2, 53.2, 52.89, 52.89, 51.98, 53.5, 53.5, 54.11, 53.5, 53.2, 
    53.5, 53.81, 54.11, 53.81, 54.11, 53.81, 54.11, 53.81, 53.81, 53.5, 
    54.11, 53.81, 53.81, 53.81, 54.42, 54.11, 53.5, 54.11, 53.81, 54.11, 
    54.11, 53.81, 48.62, 48.93, 48.62, 50.45, 51.37, 51.06, 51.06, 50.76, 
    50.76, 51.06, 51.06, 51.06, 51.98, 51.98, 51.98, 51.67, 51.98, 51.67, 
    51.37, 51.37, 51.67, 51.67, 51.67, 51.67, 51.67, 51.67, 51.06, 51.06, 
    51.06, 51.06, 51.06, 51.06, 51.37, 50.76, 51.06, 51.06, 50.76, 51.06, 
    51.06, 51.06, 50.45, 50.76, 50.45, 50.15, 49.84, 49.84, 49.84, 49.84, 
    49.23, 49.54, 49.54, 49.54, 49.84, 50.76, 51.06, 50.76, 50.76, 51.06, 
    51.06, 51.06, 51.06, 51.06, 51.06, 51.06, 51.37, 51.06, 50.76, 50.45, 
    50.45, 50.45, 50.45, 50.15, 50.15, 49.54, 49.23, 48.32, 47.71, 47.71, 
    47.4, 47.4, 47.71, 50.45, 51.06, 50.76, 51.06, 51.06, 50.76, 51.06, 
    51.06, 50.45, 50.76, 51.06, 50.76, 51.06, 51.06, 51.06, 50.76, 51.06, 
    50.76, 51.06, 50.76, 54.42, 53.81, 54.42, 55.03, 54.72, 54.72, 54.72, 
    54.11, 54.11, 53.81, 54.72, 54.11, 54.72, 54.42, 54.11, 54.11, 54.72, 
    53.81, 53.81, 54.42, 54.72, 54.42, 55.03, 54.42, 55.03, 55.03, 54.72, 
    54.72, 53.81, 54.72, 55.03, 54.72, 54.72, 54.42, 54.11, 54.72, 54.11, 
    54.72, 54.42, 54.42, 54.72, 54.72, 54.42, 54.72, 55.03, 55.03, 55.03, 
    54.72, 54.42, 54.72, 54.72, 53.81, 54.11, 54.72, 55.03, 54.72, 54.72, 
    53.81, 54.42, 54.72, 54.11, 55.03, 55.03, 55.03, 55.03, 54.11, 53.5, 
    55.03, 55.03, 54.72, 55.03, 54.72, 54.11, 54.72, 55.03, 54.72, 54.42, 
    54.72, 54.72, 55.03, 54.42, 54.11, 53.81, 53.81, 54.72, 54.11, 55.03, 
    54.42, 54.42, 53.81, 55.03, 55.03, 54.72, 54.72, 54.72, 54.42, 54.72, 
    54.72, 54.11, 54.11, 53.81, 53.81, 53.81, 53.81, 54.72, 52.89, 53.2, 
    52.59, 53.2, 52.59, 52.89, 53.2, 51.98, 51.67, 51.98, 51.37, 52.28, 
    51.98, 51.98, 52.28, 52.28, 52.28, 51.98, 51.98, 52.28, 51.98, 52.28, 
    51.67, 51.67, 51.67, 52.59, 52.28, 51.67, 51.67, 51.98, 51.98, 51.67, 
    51.37, 49.84, 48.32, 53.5, 53.2, 53.2, 52.89, 53.2, 52.89, 52.89, 52.89, 
    52.59, 52.28, 52.28, 52.59, 52.59, 52.89, 52.59, 52.59, 52.59, 52.59, 
    52.28, 52.28, 51.98, 52.59, 52.28, 52.28, 52.28, 52.28, 52.28, 51.98, 
    52.28, 52.28, 51.98, 51.98, 52.59, 51.98, 52.28, 51.98, 52.59, 51.98, 
    51.98, 51.98, 51.98, 51.67, 52.28, 51.67, 51.98, 51.98, 51.67, 51.98, 
    51.98, 51.67, 51.98, 51.67, 51.67, 51.98, 51.67, 51.98, 51.98, 51.98, 
    51.37, 51.67, 51.06, 51.67, 51.67, 51.37, 51.67, 51.67, 53.5, 54.72, 
    55.34, 55.03, 55.34, 55.34, 54.72, 55.03, 54.42, 55.34, 55.03, 54.11, 
    54.72, 54.11, 54.42, 54.42, 54.42, 54.42, 55.03, 54.72, 55.03, 53.81, 
    54.72, 54.42, 55.03, 54.72, 54.11, 53.81, 54.72, 54.72, 54.11, 54.72, 
    54.42, 54.42, 53.81, 54.42, 54.11, 54.11, 54.42, 53.81, 53.81, 54.11, 
    54.42, 54.42, 53.2, 54.42, 53.81, 54.42, 54.42, 53.81, 54.42, 54.11, 
    54.11, 54.11, 54.42, 54.42, 54.11, 55.64, 55.34, 55.34, 54.72, 55.64, 
    55.64, 55.03, 54.42, 55.34, 55.64, 55.64, 54.42, 55.34, 55.64, 55.95, 
    55.64, 55.03, 55.34, 55.64, 55.34, 55.34, 55.03, 54.42, 54.72, 54.72, 
    55.03, 54.42, 55.03, 54.42, 55.34, 55.03, 55.03, 55.34, 53.81, 55.34, 
    55.34, 55.03, 55.03, 55.03, 55.34, 55.03, 54.42, 54.72, 54.72, 54.72, 
    54.42, 55.34, 55.03, 55.34, 55.03, 55.03, 55.03, 54.72, 54.72, 54.42, 
    55.03, 55.03, 54.72, 55.03, 55.03, 54.72, 55.34, 55.03, 54.72, 54.72, 
    55.03, 54.72, 54.72, 54.11, 54.72, 54.42, 53.81, 54.72, 53.5, 53.81, 
    53.81, 54.42, 54.42, 54.42, 53.81, 54.72, 54.72, 54.72, 54.42, 54.42, 
    54.11, 54.11, 54.11, 53.5, 54.11, 54.72, 53.81, 53.81, 54.11, 53.81, 
    54.72, 54.42, 54.11, 54.72, 54.42, 54.42, 53.81, 54.42, 54.72, 54.42, 
    53.81, 53.81, 54.42, 54.42, 54.11, 54.72, 53.2, 53.2, 54.11, 54.11, 
    54.42, 54.11, 54.42, 54.11, 54.11, 53.5, 53.81, 54.42, 53.5, 54.11, 
    54.42, 53.5, 54.42, 54.42, 54.11, 53.81, 54.11, 54.42, 54.11, 54.11, 
    54.11, 54.11, 54.42, 54.11, 53.5, 54.42, 54.42, 54.11, 54.11, 53.5, 
    54.11, 53.81, 54.42, 54.11, 54.42, 54.11, 53.81, 54.11, 54.11, 54.11, 
    54.11, 54.11, 53.81, 53.2, 53.81, 52.89, 53.2, 53.5, 53.5, 53.5, 53.81, 
    53.81, 54.11, 53.81, 53.81, 54.11, 53.81, 53.81, 54.11, 53.81, 53.81, 
    53.81, 53.81, 53.81, 53.5, 53.81, 53.2, 53.2, 53.5, 53.5, 53.81, 53.81, 
    53.2, 53.81, 53.2, 53.2, 53.81, 53.2, 53.5, 54.11, 54.11, 54.11, 54.11, 
    53.5, 52.89, 53.81, 54.11, 53.81, 53.81, 53.5, 53.2, 52.89, 52.89, 53.81, 
    54.11, 54.11, 54.11, 53.5, 53.81, 54.11, 54.11, 53.81, 53.2, 53.2, 53.2, 
    53.81, 53.81, 53.81, 52.89, 53.2, 53.81, 53.2, 53.2, 52.89, 53.5, 53.5, 
    53.81, 53.81, 52.89, 54.11, 53.5, 53.81, 53.5, 53.81, 51.67, 51.37, 
    51.37, 51.67, 51.37, 51.06, 51.37, 51.06, 51.06, 51.06, 51.37, 51.06, 
    51.37, 54.42, 55.03, 54.72, 54.11, 54.72, 54.42, 54.72, 55.03, 55.03, 
    54.11, 55.03, 55.03, 53.81, 54.11, 54.72, 54.72, 55.03, 54.72, 53.81, 
    54.72, 54.72, 54.72, 53.81, 55.03, 54.42, 55.03, 54.72, 54.72, 55.03, 
    55.03, 54.72, 54.72, 54.72, 54.72, 54.72, 54.42, 54.42, 54.42, 53.5, 
    54.72, 54.11, 53.81, 54.72, 53.81, 53.5, 54.42, 54.72, 54.11, 54.42, 
    55.03, 54.11, 54.42, 54.11, 54.72, 54.72, 53.5, 53.5, 54.72, 55.03, 
    55.03, 54.72, 55.03, 54.42, 54.72, 54.42, 54.72, 55.03, 54.72, 54.72, 
    55.03, 54.11, 54.11, 54.72, 54.72, 55.03, 54.72, 55.03, 54.72, 54.72, 
    54.42, 54.42, 54.42, 54.11, 54.11, 53.81, 55.03, 53.81, 54.11, 54.72, 
    54.72, 54.72, 55.03, 55.03, 54.72, 54.72, 54.72, 54.72, 54.72, 55.03, 
    55.03, 54.72, 54.11, 54.72, 53.81, 54.11, 55.03, 54.72, 54.42, 55.03, 
    54.72, 55.03, 55.03, 54.72, 54.72, 55.03, 54.72, 54.42, 55.03, 54.42, 
    54.42, 54.72, 54.72, 54.72, 54.42, 54.42, 54.11, 54.72, 54.11, 54.72, 
    54.72, 53.81, 54.11, 54.42, 54.42, 54.72, 54.72, 54.42, 53.81, 54.42, 
    54.72, 53.5, 54.42, 54.72, 54.72, 54.72, 54.72, 54.72, 54.42, 50.76, 
    50.76, 50.76, 50.76, 50.76, 51.06, 51.06, 50.76, 50.76, 50.45, 50.45, 
    50.15, 50.45, 50.45, 51.06, 51.06, 51.06, 50.76, 51.06, 50.76, 50.76, 
    50.76, 50.15, 50.45, 50.45, 50.45, 50.45, 50.76, 49.84, 49.84, 49.84, 
    50.15, 49.84, 49.84, 49.84, 49.54, 49.84, 49.54, 49.54, 49.23, 49.54, 
    49.54, 49.84, 49.84, 49.84, 49.84, 49.84, 49.54, 49.54, 49.23, 49.54, 
    49.84, 49.54, 52.59, 55.34, 55.03, 55.34, 54.42, 55.34 ;

 IP = 0, 8.64, 5.9, 0.4, 0, 0, 0, 0, 0, 0, 0, 23.29, 24.82, 10.47, 25.73, 
    21.46, 13.83, 13.83, 12.61, 8.03, 1.93, 2.54, 0.4, 2.54, 0, 15.97, 23.29, 
    20.24, 29.39, 22.99, 25.12, 15.66, 20.24, 12.92, 21.46, 20.85, 28.48, 
    17.8, 20.54, 25.73, 23.6, 30.62, 23.29, 16.58, 21.77, 16.27, 12.61, 
    12.61, 11.39, 10.78, 3.76, 7.42, 3.45, 7.12, 5.9, 6.81, 2.23, 0.1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.71, 6.81, 21.16, 4.68, 0.1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.01, 0, 0.4, 0.4, 0, 0.1, 0, 0, 0, 0, 
    0, 0, 0, 0, 3.76, 24.51, 2.23, 7.42, 3.15, 9.56, 12.92, 22.07, 9.56, 
    10.47, 5.29, 1.93, 0, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 1.01, 4.37, 19.63, 
    8.34, 0.4, 0, 0, 0, 0, 0, 0, 5.9, 12.61, 7.73, 22.38, 7.73, 1.32, 12.3, 
    8.34, 0.71, 0.4, 0, 0, 0, 0, 1.62, 24.82, 4.98, 0, 0, 0, 0, 0, 0, 0, 0.1, 
    0, 12.61, 26.04, 23.29, 3.45, 2.54, 0.1, 0, 0, 1.93, 2.84, 2.23, 22.68, 
    19.02, 24.21, 8.95, 23.6, 30.62, 24.82, 16.88, 19.93, 24.51, 27.56, 
    25.73, 15.05, 23.29, 24.21, 5.9, 6.81, 5.59, 6.2, 10.47, 20.85, 11.39, 
    24.82, 21.46, 27.26, 27.56, 27.56, 24.21, 19.32, 19.32, 19.63, 8.95, 
    1.32, 1.32, 5.59, 1.93, 0, 0.71, 1.93, 0, 0.71, 2.84, 8.03, 17.8, 26.04, 
    26.34, 25.12, 29.7, 24.51, 26.04, 24.82, 23.6, 25.12, 25.43, 20.24, 
    11.08, 16.27, 10.78, 13.53, 3.15, 1.01, 0, 0.4, 1.62, 25.73, 9.56, 4.37, 
    17.19, 21.46, 19.32, 26.95, 17.19, 16.58, 6.51, 7.12, 6.81, 0.1, 12.61, 
    7.73, 14.75, 20.85, 26.34, 12.3, 25.12, 7.73, 12, 20.54, 21.77, 12, 
    20.54, 8.34, 8.34, 8.95, 4.98, 12.61, 2.84, 2.84, 1.93, 0.1, 3.45, 8.34, 
    2.54, 18.41, 2.54, 28.17, 7.73, 6.81, 20.24, 22.68, 22.68, 12.92, 9.56, 
    10.78, 12, 8.95, 14.44, 3.45, 27.26, 19.93, 17.19, 14.75, 9.25, 7.42, 
    8.64, 7.73, 1.62, 5.29, 5.59, 4.07, 1.93, 0.1, 3.76, 1.01, 1.32, 1.93, 
    1.93, 1.93, 1.32, 5.29, 3.15, 1.62, 4.37, 24.21, 5.59, 13.83, 6.2, 15.05, 
    30.31, 12.3, 6.51, 19.02, 6.51, 17.49, 8.34, 12.92, 2.23, 4.07, 4.68, 
    1.62, 1.32, 8.95, 8.95, 6.2, 2.84, 3.45, 1.32, 5.9, 14.14, 7.12, 15.05, 
    3.76, 1.32, 8.34, 6.51, 3.76, 3.76, 13.22, 11.69, 1.62, 1.62, 0.71, 
    16.27, 1.93, 3.76, 1.93, 12.92, 13.83, 14.75, 26.34, 12.92, 3.76, 2.84, 
    1.32, 4.98, 8.95, 8.34, 13.83, 10.78, 13.22, 11.69, 14.14, 21.77, 21.46, 
    22.07, 21.16, 17.8, 18.41, 18.1, 9.25, 20.24, 14.75, 15.05, 9.56, 12.3, 
    26.04, 30.62, 15.97, 10.47, 25.43, 16.27, 18.1, 21.16, 12.92, 21.46, 
    28.48, 20.54, 19.93, 23.9, 19.63, 21.16, 22.07, 15.97, 16.88, 18.71, 
    11.39, 12.61, 6.2, 7.12, 8.95, 6.51, 6.81, 3.76, 4.68, 4.98, 1.93, 1.32, 
    3.76, 18.1, 11.69, 13.83, 19.93, 11.08, 11.39, 16.27, 13.53, 19.32, 
    14.44, 14.75, 24.21, 17.8, 20.24, 13.53, 18.1, 21.46, 26.65, 16.58, 
    15.97, 11.39, 18.71, 6.2, 8.95, 7.42, 12.61, 10.78, 7.73, 5.9, 7.42, 
    7.42, 7.12, 8.03, 7.73, 10.78, 9.86, 10.78, 6.51, 11.39, 7.42, 6.81, 6.2, 
    2.54, 3.15, 4.07, 3.45, 3.45, 3.76, 4.37, 2.84, 3.76, 3.45, 3.15, 1.93, 
    2.23, 0.71, 1.01, 2.84, 0, 0.4, 0.71, 0.1, 0, 1.01, 0, 0, 0, 0.1, 0, 0.4, 
    0, 1.32, 0, 0, 0.1, 0.1, 0, 0, 0, 0, 0, 0, 0.1, 0, 0.1, 0.1, 0, 0.4, 0, 
    0, 0, 0, 0, 0, 3.76, 0.1, 1.01, 0, 0.1, 0.4, 0.4, 0, 4.98, 0, 1.01, 0.71, 
    2.23, 19.63, 22.38, 8.03, 1.32, 1.01, 0.71, 0, 0, 0, 0.71, 0, 0, 0, 0.4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.01, 0, 3.15, 0, 0, 1.01, 0, 0, 0.1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.07, 6.2, 19.93, 13.83, 
    12.61, 4.07, 1.62, 0.4, 8.95, 2.54, 1.62, 4.07, 7.42, 6.51, 3.76, 2.54, 
    5.9, 5.29, 7.12, 3.76, 4.07, 2.23, 2.23, 17.8, 3.15, 5.29, 11.39, 1.62, 
    1.01, 0.4, 0, 0.1, 0.1, 0, 0, 0, 0.4, 0.1, 0, 0.71, 0, 0.4, 0.71, 0.1, 
    0.4, 4.98, 22.68, 19.32, 9.86, 25.43, 28.78, 22.38, 28.48, 37.02, 14.44, 
    26.95, 19.93, 11.69, 14.14, 11.08, 11.08, 14.44, 8.03, 8.03, 3.76, 8.64, 
    4.68, 1.93, 1.01, 0.4, 0.4, 0.1, 0, 0, 0, 0, 0.1, 0.1, 1.62, 16.27, 
    10.47, 23.6, 17.49, 5.29, 0.1, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0.1, 
    0, 1.62, 1.01, 18.41, 24.51, 4.98, 2.23, 0.1, 0, 0.4, 0.1, 2.54, 0, 0.1, 
    0, 0, 0, 0, 0, 0, 0.1, 0.1, 0.4, 4.07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.01, 2.23, 15.66, 2.54, 3.15, 3.76, 1.32, 5.59, 3.15, 2.54, 2.23, 8.64, 
    15.36, 11.08, 2.23, 15.66, 29.09, 12.61, 12.61, 22.68, 11.08, 2.23, 1.93, 
    2.54, 2.23, 1.01, 0.4, 2.23, 0.4, 0.1, 0, 0.71, 0, 0, 0, 0, 0, 0, 0.1, 
    24.21, 14.14, 2.23, 0.1, 0, 1.62, 0, 0, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 0.4, 
    9.86, 6.81, 10.17, 10.17, 21.46, 10.47, 1.62, 5.29, 5.29, 9.56, 9.56, 
    12.3, 3.76, 2.54, 3.15, 0.71, 1.01, 0.4, 0.4, 0, 0, 0.1, 0, 0.4, 0, 0.71, 
    0.4, 0, 0.4, 0.71, 0.1, 1.01, 0.71, 0.1, 1.93, 1.32, 0.1, 0, 0, 0.1, 0, 
    0.4, 0, 0, 0, 0, 0, 0, 0.4, 0.71, 2.84, 14.75, 15.66, 2.54, 4.07, 7.42, 
    8.64, 1.01, 1.93, 2.84, 5.9, 5.9, 23.29, 18.71, 8.95, 11.69, 11.69, 6.2, 
    3.45, 7.12, 0.4, 0.4, 0.1, 0, 0.4, 0.71, 0.4, 0, 0.4, 0.4, 0.1, 0.4, 
    1.32, 4.07, 4.68, 0, 0.4, 0, 0.1, 0.1, 0, 0, 0, 0, 0.1, 0.1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0.1, 0, 0, 0, 0, 0, 
    0, 0, 0.1, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0.71, 0.71, 0.4, 
    0.1, 0.4, 0.4, 6.81, 3.76, 6.2, 2.54, 1.01, 0.4, 1.32, 0, 0, 0, 0.1, 0, 
    0.4, 0.1, 0, 0, 0, 0, 0, 16.58, 19.02, 1.32, 0.1, 0.1, 0.4, 0.1, 0, 0, 
    0.1, 1.93, 10.78, 9.56, 0.4, 1.01, 0.71, 3.76, 5.9, 15.36, 3.45, 22.07, 
    4.68, 1.62, 0, 0, 0, 0, 0, 0, 0, 0, 13.83, 0.1, 0, 0.1, 0, 0, 0.1, 0, 0, 
    7.42, 2.23, 0.4, 0.4, 0, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 
    0.1, 0.1, 0.71, 0, 2.23, 1.32, 0.1, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.4, 0.71, 1.01, 0.71, 0, 0, 0, 0.1, 0.4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7.12, 0, 0, 1.62, 2.23, 15.97, 0, 0.1, 0, 0, 0.4, 16.88, 0.71, 0.1, 
    0, 0, 0, 0, 0, 0.1, 0, 0, 4.37, 11.69, 0.4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0.1, 0, 0, 0, 0, 0, 0, 1.01, 0, 0, 0, 0.1, 
    0, 0, 0, 0, 0.1, 0, 1.01, 2.54, 0, 0.1, 0.4, 0, 0, 0, 0, 0, 0, 1.32, 
    8.34, 10.47, 1.62, 0.4, 1.01, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.71, 0.1, 0.71, 0, 0, 0.1, 0, 0.1, 0, 0.1, 0, 0, 0.1, 0.4, 0, 21.46, 
    4.07, 0.71, 1.32, 0.1, 0, 0.1, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0.1, 
    1.32, 2.84, 0.1, 0, 0, 0, 0, 0, 0.1, 0, 0.71, 9.86, 0.71, 0.4, 0, 0, 0, 
    0, 0, 0.1, 0, 0, 0.1, 0, 0, 0, 0, 0.4, 0.4, 14.44, 0.1, 0.1, 0.4, 0.1, 0, 
    0.1, 0, 0, 4.07, 8.34, 2.23, 4.37, 3.15, 8.03, 0.1, 0, 0.1, 0 ;

 TQ = 41.6, 30.01, 32.45, 20.85, 20.85, 25.43, 20.85, 21.77, 24.82, 21.77, 
    30.92, 33.67, 30.31, 20.24, 26.34, 28.48, 30.92, 33.97, 30.62, 35.8, 
    24.82, 26.65, 27.26, 25.12, 29.39, 35.8, 32.14, 32.75, 25.12, 22.38, 
    28.17, 22.68, 26.04, 26.95, 29.39, 30.62, 32.14, 24.21, 30.92, 27.26, 
    25.12, 32.14, 27.26, 26.95, 27.87, 26.34, 28.17, 29.09, 24.51, 26.04, 
    28.48, 24.51, 33.97, 31.53, 30.92, 28.78, 22.99, 21.77, 19.02, 19.93, 
    8.03, 18.1, 14.44, 22.68, 16.88, 13.83, 19.93, 18.41, 30.62, 36.11, 
    34.89, 36.41, 35.5, 26.65, 33.67, 41.3, 19.32, 32.45, 54.42, 17.49, 18.1, 
    12, 29.39, 30.62, 21.77, 23.9, 24.51, 25.12, 31.84, 25.43, 28.78, 32.75, 
    34.28, 33.36, 28.78, 29.09, 28.48, 27.26, 31.23, 21.77, 37.94, 27.26, 
    26.34, 30.31, 29.39, 34.89, 30.01, 33.36, 34.89, 32.75, 35.19, 33.36, 
    35.19, 31.53, 27.26, 21.46, 43.43, 37.33, 22.38, 9.86, 33.67, 8.03, 
    36.41, 29.39, 17.49, 24.82, 28.17, 34.28, 33.67, 37.02, 31.84, 21.16, 
    32.75, 21.77, 28.48, 33.06, 26.65, 32.75, 38.86, 39.16, 31.84, 38.25, 
    33.36, 35.8, 41.6, 33.97, 24.21, 40.08, 26.65, 36.72, 32.14, 38.25, 
    43.43, 37.94, 26.65, 27.87, 20.24, 15.36, 25.12, 24.82, 22.38, 29.09, 
    33.67, 29.7, 38.55, 41.91, 27.26, 32.14, 30.92, 33.06, 26.04, 25.73, 
    28.17, 28.78, 33.36, 37.94, 39.16, 35.19, 33.67, 31.84, 26.65, 35.5, 
    29.7, 29.39, 31.23, 36.72, 36.72, 25.12, 30.01, 25.73, 36.41, 43.13, 
    34.28, 38.55, 36.11, 34.89, 30.62, 29.09, 33.06, 29.39, 26.65, 26.04, 
    31.84, 26.65, 27.87, 20.24, 31.84, 33.67, 26.34, 40.99, 35.8, 39.47, 
    29.7, 33.67, 36.41, 42.21, 40.69, 30.62, 30.31, 23.6, 26.34, 25.43, 23.9, 
    26.95, 32.14, 37.33, 28.48, 24.21, 30.92, 29.39, 38.86, 33.67, 33.97, 
    41.6, 31.53, 33.36, 30.01, 35.8, 33.06, 31.53, 32.45, 32.75, 33.67, 
    34.28, 26.95, 26.95, 30.01, 32.45, 32.45, 30.92, 28.78, 29.09, 34.28, 
    34.28, 32.45, 26.95, 29.39, 33.97, 26.65, 30.92, 31.53, 30.01, 27.26, 
    30.01, 38.55, 30.62, 35.8, 37.94, 34.58, 35.5, 31.84, 29.7, 30.31, 32.75, 
    28.48, 33.06, 29.09, 31.53, 26.34, 27.26, 35.19, 39.77, 33.06, 26.95, 
    28.78, 26.04, 28.17, 26.65, 23.6, 26.95, 27.87, 30.62, 24.51, 31.23, 
    31.53, 26.34, 34.28, 30.62, 28.17, 30.92, 28.78, 30.62, 29.7, 35.19, 
    28.17, 30.01, 24.51, 28.78, 30.62, 30.31, 25.12, 29.39, 30.92, 27.87, 
    30.31, 27.26, 26.34, 26.65, 30.92, 31.23, 31.53, 31.23, 22.99, 28.78, 
    33.06, 30.62, 36.72, 28.17, 33.67, 33.36, 38.25, 32.75, 24.82, 27.56, 
    37.02, 32.45, 33.36, 27.56, 30.92, 27.26, 33.67, 31.84, 30.31, 26.95, 
    31.53, 30.92, 34.58, 33.67, 29.09, 30.92, 24.82, 32.75, 31.53, 31.53, 
    27.56, 28.78, 27.87, 26.65, 30.31, 28.17, 25.43, 28.17, 35.8, 31.23, 
    26.04, 39.16, 31.53, 37.94, 38.55, 36.72, 44.04, 35.19, 39.47, 38.25, 
    35.8, 35.19, 38.86, 37.94, 44.35, 77.31, 27.56, 24.21, 23.29, 27.87, 
    25.73, 33.06, 28.17, 33.36, 29.09, 31.23, 30.62, 27.56, 33.67, 30.31, 
    28.78, 28.48, 35.5, 26.95, 31.84, 32.75, 25.73, 25.73, 34.28, 27.56, 
    27.56, 21.77, 29.09, 29.39, 25.12, 30.01, 30.92, 30.01, 29.39, 30.62, 
    33.36, 28.17, 27.87, 24.82, 25.43, 25.43, 33.67, 34.89, 36.11, 34.28, 
    28.17, 28.17, 30.01, 28.78, 28.78, 28.78, 33.06, 37.94, 36.41, 34.58, 
    21.16, 26.04, 26.95, 28.17, 32.45, 22.99, 22.38, 29.39, 28.78, 33.06, 
    37.94, 32.14, 25.43, 25.73, 25.73, 26.95, 29.39, 32.14, 28.17, 29.7, 
    28.48, 27.26, 24.51, 22.38, 21.77, 22.07, 21.77, 32.75, 31.84, 26.34, 
    41.91, 26.65, 33.36, 44.65, 43.43, 40.69, 36.11, 48.32, 44.65, 45.57, 
    43.43, 43.74, 33.36, 34.28, 35.19, 36.72, 19.93, 19.32, 20.54, 27.87, 
    41.3, 25.43, 50.76, 29.09, 8.64, 17.8, 24.51, 33.67, 32.14, 62.35, 24.21, 
    33.97, 43.43, 46.49, 26.04, 28.17, 46.79, 28.48, 36.11, 37.02, 27.56, 
    25.12, 24.51, 35.8, 40.38, 39.47, 22.38, 26.95, 16.88, 33.67, 22.99, 
    27.26, 29.7, 33.97, 31.23, 31.23, 27.87, 30.31, 26.04, 34.89, 33.67, 
    27.87, 26.95, 29.7, 29.39, 42.21, 38.86, 31.23, 39.47, 34.58, 26.65, 
    42.52, 25.73, 35.5, 33.36, 28.78, 30.31, 37.33, 40.38, 30.92, 26.65, 
    27.56, 29.7, 24.82, 31.84, 28.17, 23.9, 27.56, 26.34, 30.62, 37.63, 
    36.41, 26.65, 27.87, 22.99, 31.23, 22.38, 22.68, 21.16, 17.49, 21.77, 
    26.95, 17.19, 20.85, 33.97, 10.78, 14.44, 25.43, 20.24, 27.87, 37.02, 
    33.36, 24.51, 19.63, 30.31, 39.16, 36.72, 35.19, 35.8, 30.92, 37.33, 
    41.3, 42.82, 38.86, 42.82, 51.98, 53.2, 38.86, 44.04, 56.25, 45.87, 
    40.69, 33.67, 33.06, 37.33, 45.57, 41.91, 44.96, 45.26, 33.06, 38.55, 
    33.97, 40.38, 27.87, 29.39, 48.01, 29.09, 33.97, 24.82, 26.95, 23.9, 
    27.26, 33.36, 25.12, 25.43, 25.43, 25.12, 31.53, 27.87, 25.12, 28.78, 
    29.7, 26.95, 22.99, 28.78, 31.84, 27.87, 28.48, 22.68, 24.21, 33.67, 
    32.14, 27.87, 28.48, 33.06, 34.28, 34.89, 44.65, 37.02, 32.45, 37.33, 
    38.86, 29.39, 29.7, 25.73, 28.48, 30.31, 32.45, 36.41, 39.16, 35.5, 
    33.97, 32.45, 33.97, 35.5, 36.72, 43.74, 42.52, 43.74, 34.58, 34.58, 
    25.12, 33.97, 36.41, 34.58, 29.7, 33.67, 42.82, 41.91, 36.41, 30.92, 
    38.25, 26.95, 30.31, 35.5, 33.67, 36.41, 35.8, 34.58, 33.36, 35.8, 30.62, 
    29.09, 29.7, 28.17, 34.28, 32.75, 35.19, 29.39, 29.39, 32.14, 26.95, 
    38.86, 42.52, 33.06, 33.36, 35.5, 30.01, 28.78, 34.58, 35.19, 30.01, 
    28.78, 26.95, 27.56, 19.32, 18.1, 22.07, 31.84, 34.89, 28.78, 29.7, 
    30.31, 26.95, 30.31, 30.92, 31.23, 30.92, 28.48, 31.53, 32.75, 33.97, 
    32.75, 32.45, 32.75, 33.06, 42.82, 37.94, 36.72, 38.55, 36.41, 26.34, 
    29.39, 26.95, 29.7, 29.09, 28.17, 30.62, 24.82, 34.89, 27.56, 28.78, 
    24.51, 29.09, 27.56, 30.31, 28.78, 44.35, 34.58, 28.17, 32.75, 29.09, 
    29.39, 26.34, 24.21, 28.78, 27.26, 27.56, 23.29, 22.68, 40.38, 32.45, 
    34.58, 30.01, 33.67, 38.55, 34.28, 32.45, 32.45, 37.02, 37.94, 35.8, 
    39.47, 37.02, 39.47, 36.72, 32.14, 26.04, 29.39, 30.31, 28.48, 24.51, 
    27.87, 28.78, 25.12, 22.07, 27.56, 27.56, 24.21, 25.12, 25.12, 25.73, 
    25.12, 30.62, 32.14, 29.39, 28.17, 27.87, 28.17, 22.38, 24.21, 19.32, 
    24.21, 25.12, 24.82, 30.62, 23.29, 26.04, 28.17, 26.65, 25.12, 22.99, 
    29.39, 33.97, 31.53, 36.11, 32.75, 29.09, 32.14, 41.6, 38.86, 32.14, 
    38.55, 42.82, 42.21, 37.63, 34.89, 44.96, 32.45, 36.41, 34.89, 32.45, 
    28.17, 28.17, 28.78, 31.53, 23.9, 23.9, 26.65, 27.26, 28.48, 27.87, 
    25.12, 25.43, 30.01, 29.09, 28.17, 28.17, 22.07, 26.95, 27.26, 28.78, 
    31.53, 30.31, 23.9, 26.65, 29.09, 23.9, 42.21, 23.29, 30.31, 33.97, 
    26.34, 35.8, 25.73, 22.07, 41.6, 41.3, 25.73, 15.97, 30.31, 26.95, 30.01, 
    22.99, 34.28, 33.67, 19.32, 19.02, 18.1, 23.9, 18.41, 20.54, 20.85, 
    21.46, 21.77, 21.77, 34.28, 27.26, 26.34, 18.71, 20.85, 23.29, 18.71, 
    15.66, 21.46, 28.48, 19.02, 20.54, 21.46, 28.78, 36.41, 43.13, 25.12, 
    17.49, 36.41, 22.99, 51.37, 51.06, 49.54, 34.28, 36.41, 28.78, 26.04, 
    37.33, 39.16, 28.17, 27.56, 37.33, 40.69, 60.22, 21.77, 19.93, 22.38, 
    19.02, 25.73, 30.01, 41.6, 36.41, 30.31, 45.26, 23.9, 18.41, 25.12, 
    25.73, 21.77, 20.85, 31.53, 38.55, 38.55, 22.99, 32.75, 31.53, 52.59, 
    37.63, 38.25, 40.38, 41.6, 37.02, 45.57, 19.93, 30.01, 30.31, 21.16, 
    22.38, 20.54, 26.34, 29.09, 35.19, 44.65, 21.77, 29.7, 27.56, 23.29, 
    30.31, 23.9, 27.87, 34.89, 44.65, 33.06, 32.45, 33.36, 41.6, 39.77, 
    32.14, 20.54, 23.9, 25.73, 21.77, 23.9, 18.41, 19.93, 15.05, 24.82, 23.9, 
    22.07, 36.72, 26.04, 27.56, 30.01, 35.5, 35.5, 33.36, 40.38, 21.16, 
    33.06, 24.21, 34.89, 25.43, 35.19, 19.02, 27.56, 33.67, 37.94, 45.26, 
    34.89, 34.89, 31.84, 19.93, 22.38, 26.34, 27.87, 38.86, 33.36, 37.94, 
    28.78, 18.1, 30.92, 21.46, 26.04, 21.77, 25.12, 22.07, 20.24, 40.08, 
    44.35, 39.16, 18.71, 23.9, 30.62, 50.15, 23.29, 20.24, 33.67, 30.01, 
    33.67, 49.84, 31.84, 29.09, 28.78, 30.62, 22.99, 25.12, 24.82, 26.65, 
    27.87, 32.45, 35.8, 38.25, 38.25, 51.98, 32.75, 38.55, 40.99, 32.14, 
    34.28, 23.6, 29.39, 32.14, 34.28, 43.74, 39.77, 33.36, 32.14, 24.82, 
    47.1, 32.45, 35.8, 26.65, 31.84, 30.62, 46.18, 27.26, 27.26, 34.28, 
    40.38, 52.28, 21.46, 40.38, 32.45, 35.5, 36.72, 43.13, 27.87, 25.73, 
    34.89, 32.45, 41.6, 47.4, 35.8, 23.29, 29.09, 28.48, 29.7, 21.46, 27.87, 
    29.7, 37.02, 41.91, 47.4, 40.38, 40.69, 33.36, 41.6, 40.99, 54.42, 48.93, 
    28.17, 25.73, 19.32, 31.84, 38.25, 26.04, 19.63, 32.75, 40.08, 43.74, 
    38.86, 41.3, 68.46, 34.28, 38.25, 40.69, 31.53, 19.32, 26.95, 36.11, 
    29.39, 28.48, 45.26, 51.06, 41.91, 60.22, 34.58, 37.63, 31.23, 54.11, 
    36.72, 51.06, 44.96, 46.49, 12.61, 37.94, 23.9, 26.65, 22.68, 29.7, 
    24.82, 26.34, 26.04, 42.82, 70.59, 27.56, 23.6, 26.04, 20.85, 30.92, 
    32.75, 18.71, 30.92, 15.97, 35.5, 46.18, 41.3, 30.01, 59.91, 40.69, 
    30.62, 41.3, 26.04, 22.07, 30.92, 30.31, 30.31, 18.1, 21.46, 29.7, 22.99, 
    50.15, 44.35, 37.02, 33.67, 21.77, 19.93, 30.92, 28.17, 22.07, 13.22, 
    38.86, 40.69, 53.5, 37.94, 41.6, 32.14, 33.06, 33.06, 25.12, 33.97, 
    28.17, 35.19 ;

 HP = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 
    0, 0.1, 0, 0, 0.1, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0.1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 
    0, 0.1, 0, 0, 0, 0.1, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 
    0.1, 0.1, 0.1, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 0, 
    0, 0.1, 0, 0, 0.1, 0, 0, 0, 0, 0.1, 0, 0, 0.1, 0, 0, 0.1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 0.1, 0, 0.1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0.1, 0.1, 0, 0, 0, 0, 0.1, 0, 0, 
    0.1, 0, 0, 0.1, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 0.1, 0, 
    0.1, 0, 0, 0.1, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0.1, 0, 0, 0, 
    0, 0.1, 0.1, 0, 0, 0, 0.1, 0, 0, 0, 0, 0.1, 0, 0.1, 0.1, 0, 0.1, 0, 0.1, 
    0, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0, 0.1, 0, 0, 0, 0, 
    0, 0.1, 0.1, 0, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 0, 0.1, 0.1, 0.1, 0, 0.1, 0, 
    0, 0.1, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 0, 0.1, 0, 0.1, 0.1, 0, 0, 0, 0, 0.1, 
    0.1, 0, 0, 0, 0.1, 0, 0, 0, 0, 0.1, 0.1, 0.1, 0, 0, 0.1, 0, 0, 0.1, 0, 0, 
    0.1, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0, 0, 0, 0, 0.1, 0.1, 0.1, 0, 
    0.1, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 0, 
    0, 0, 0, 0, 0, 0.1, 0.1, 0, 0.1, 0, 0.1, 0.1, 0, 0.1, 0, 0.1, 0, 0.1, 
    0.1, 0.1, 0.4, 0.4, 0.4, 0.4, 0.4, 0.1, 0, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0, 0.1, 0.1, 0, 0, 0.1, 0.1, 0, 0, 0.1, 0.1, 0.1, 0, 0.1, 0, 0, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0, 0.1, 0, 0, 0.1, 0, 0, 0.1, 0.1, 0, 0.1, 0.1, 0.1, 
    0, 0.1, 0.1, 0, 0, 0, 0, 0.1, 0.1, 0, 0, 0.1, 0.1, 0.1, 0, 0.1, 0.1, 0, 
    0, 0.1, 0.1, 0.1, 0, 0, 0.1, 0.1, 0, 0.1, 0.1, 0.1, 0, 0, 0, 0, 0.1, 0.1, 
    0, 0.1, 0, 0, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 0, 0, 0, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0, 0, 0, 0.1, 0.1, 0.1, 0.1, 0.1, 0, 0.1, 0, 0, 0.1, 0.1, 0, 0, 0.1, 
    0.1, 0.1, 0, 0, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0, 0, 0.1, 0, 0.1, 0, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 0, 0.1, 0.1, 
    0, 0.1, 0, 0.1, 0, 0.1, 0, 0.1, 0, 0, 0.1, 0.1, 0.1, 0, 0, 0, 0, 0.1, 
    0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0.1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 
    0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.1, 0.1, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 0, 0, 0.1, 0.1, 0, 0.1, 0, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0, 0, 0.1, 0, 0.1, 0, 0.1, 0.1, 0, 0, 0.1, 0.1, 0, 
    0.1, 0, 0, 0.1, 0, 0, 0, 0, 0.1, 0.1, 0, 0.1, 0, 0, 0, 0, 0, 0.1, 0, 0.1, 
    0.1, 0, 0, 0, 0, 0, 0.1, 0, 0, 0.1, 0, 0, 0, 0, 0, 0.1, 0.1, 0.1, 0, 0.1, 
    0, 0.1, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 0.1, 0.1, 0, 0, 0.1, 0, 0.1, 0.1, 
    0.1, 0, 0, 0, 0.1, 0.1, 0.1, 0.1, 0, 0.1, 0.1, 0, 0, 0, 0, 0, 0.1, 0, 
    0.1, 0, 0.1, 0, 0, 0, 0, 0, 0, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 0.1, 0, 0.1, 
    0.1, 0.1, 0, 0.1, 0, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 0.1, 0, 0, 0, 0.1, 0.1, 
    0, 0, 0.1, 0, 0.1, 0, 0, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 0, 0.1, 0, 0, 0, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
    0.4, 0.1, 0.1, 1.01, 0, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 2.23, 0.1, 0, 0, 0, 
    0.1, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0, 0.1, 0.1, 0, 
    0.1, 0, 0.1, 0, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0, 0.4, 0.4, 0.1, 
    0.1, 0, 0.1, 0.1, 0.1, 0.1, 0.1, 0, 0, 0.1, 0.1, 0.1, 0.4, 0.1, 0.1, 0.1, 
    0, 0.1, 0.1, 0.1, 0, 0.1, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 0, 0.1, 0, 0.1, 0, 
    0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0 ;
}
