netcdf data {
dimensions:
	time = UNLIMITED ; // (14 currently)
variables:
	float time(time) ;
		time:unit = "s" ;
		time:label = "time" ;
	int STEP(time) ;
		STEP:label = "Palier" ;
	float PR1(time) ;
		PR1:unit = "bar" ;
		PR1:label = "PR1S" ;
	float PR15(time) ;
		PR15:unit = "bar" ;
		PR15:label = "PR15S" ;
	float PR30(time) ;
		PR30:unit = "bar" ;
		PR30:label = "PR30S" ;
	float PR60(time) ;
		PR60:unit = "bar" ;
		PR60:label = "PR60S" ;
	float PG1(time) ;
		PG1:unit = "bar" ;
		PG1:label = "PG1S" ;
	float PG15(time) ;
		PG15:unit = "bar" ;
		PG15:label = "PG15S" ;
	float PG30(time) ;
		PG30:unit = "bar" ;
		PG30:label = "PG30S" ;
	float PG60(time) ;
		PG60:unit = "bar" ;
		PG60:label = "PG60S" ;
	float V1(time) ;
		V1:unit = "cm3" ;
		V1:label = "V1S" ;
	float V15(time) ;
		V15:unit = "cm3" ;
		V15:label = "V15S" ;
	float V30(time) ;
		V30:unit = "cm3" ;
		V30:label = "V30S" ;
	float V60(time) ;
		V60:unit = "cm3" ;
		V60:label = "V60S" ;
		V60:scale_max = 500.f ;
	float CREEP(time) ;
		CREEP:unit = "cm3" ;
		CREEP:label = "fluage" ;
	float DELT60(time) ;
		DELT60:unit = "cm3" ;
		DELT60:label = "delt60" ;
data:

 time = 80, 142, 205, 268, 330, 394, 456, 519, 582, 647, 711, 776, 840, 905 ;

 STEP = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14 ;

 PR1 = 0.06, 1.08, 1.81, 2.85, 4.01, 5.98, 7.96, 9.8, 13.87, 17.81, 22.05, 
    25.77, 29.73, 33.8 ;

 PR15 = 0.06, 0.81, 1.81, 2.82, 3.86, 5.81, 7.82, 9.81, 13.82, 17.85, 21.75, 
    25.75, 29.75, 33.76 ;

 PR30 = 0.03, 0.81, 1.82, 2.83, 3.84, 5.85, 7.82, 9.83, 13.82, 17.84, 21.78, 
    25.75, 29.77, 33.75 ;

 PR60 = 0.04, 0.82, 1.82, 2.84, 3.86, 5.83, 7.83, 9.82, 13.84, 17.81, 21.76, 
    25.75, 29.77, 33.75 ;

 PG1 = 0.11, 0.28, 1.31, 2.14, 3.17, 5.24, 7.14, 9.17, 13.21, 17.14, 21.14, 
    25.15, 29.12, 33.09 ;

 PG15 = 0.1, 0.29, 1.18, 2.12, 3.15, 5.19, 7.18, 9.17, 13.15, 17.16, 21.06, 
    25.09, 29.06, 33.08 ;

 PG30 = 0.09, 0.28, 1.19, 2.16, 3.17, 5.22, 7.17, 9.16, 13.14, 17.15, 21.1, 
    25.08, 29.1, 33.06 ;

 PG60 = 0.08, 0.29, 1.17, 2.14, 3.17, 5.18, 7.18, 9.14, 13.15, 17.13, 21.09, 
    25.08, 29.06, 33.08 ;

 V1 = 60, 103, 215, 257, 280, 303, 320, 335, 359, 386, 411, 441, 477, 518 ;

 V15 = 76, 149, 238, 266, 285, 307, 324, 339, 366, 392, 419, 452, 491, 532 ;

 V30 = 85, 176, 241, 268, 287, 308, 325, 340, 368, 395, 423, 457, 498, 540 ;

 V60 = 92, 198, 244, 270, 287, 309, 326, 342, 370, 397, 428, 463, 506, 550 ;

 CREEP = 7, 22, 3, 2, 0, 1, 1, 2, 2, 2, 5, 6, 8, 10 ;

 DELT60 = 92, 106, 46, 26, 17, 22, 17, 16, 28, 27, 31, 35, 43, 44 ;
}
