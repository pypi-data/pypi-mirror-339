netcdf data {
dimensions:
	time = UNLIMITED ; // (14 currently)
variables:
	float time(time) ;
		time:unit = "s" ;
		time:label = "time" ;
	int STEP(time) ;
		STEP:label = "Palier" ;
	float PR1(time) ;
		PR1:unit = "bar" ;
		PR1:label = "PR1S" ;
	float PR15(time) ;
		PR15:unit = "bar" ;
		PR15:label = "PR15S" ;
	float PR30(time) ;
		PR30:unit = "bar" ;
		PR30:label = "PR30S" ;
	float PR60(time) ;
		PR60:unit = "bar" ;
		PR60:label = "PR60S" ;
	float PG1(time) ;
		PG1:unit = "bar" ;
		PG1:label = "PG1S" ;
	float PG15(time) ;
		PG15:unit = "bar" ;
		PG15:label = "PG15S" ;
	float PG30(time) ;
		PG30:unit = "bar" ;
		PG30:label = "PG30S" ;
	float PG60(time) ;
		PG60:unit = "bar" ;
		PG60:label = "PG60S" ;
	float V1(time) ;
		V1:unit = "cm3" ;
		V1:label = "V1S" ;
	float V15(time) ;
		V15:unit = "cm3" ;
		V15:label = "V15S" ;
	float V30(time) ;
		V30:unit = "cm3" ;
		V30:label = "V30S" ;
	float V60(time) ;
		V60:unit = "cm3" ;
		V60:label = "V60S" ;
		V60:scale_max = 500.f ;
	float CREEP(time) ;
		CREEP:unit = "cm3" ;
		CREEP:label = "fluage" ;
	float DELT60(time) ;
		DELT60:unit = "cm3" ;
		DELT60:label = "delt60" ;
data:

 time = 78, 143, 211, 278, 348, 418, 486, 553, 622, 690, 758, 826, 897, 967 ;

 STEP = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14 ;

 PR1 = 1.09, 1.98, 3.03, 4.05, 8.59, 13.13, 17.96, 22.37, 27.2, 31.56, 36.4, 
    40.84, 45.44, 50.03 ;

 PR15 = 1.02, 1.98, 3, 3.99, 8.56, 13.16, 17.84, 22.43, 27.03, 31.56, 36.15, 
    40.77, 45.37, 50.04 ;

 PR30 = 1, 2.05, 3, 3.99, 8.55, 13.19, 17.79, 22.34, 27.03, 31.53, 36.19, 
    40.83, 45.37, 49.97 ;

 PR60 = 1, 1.94, 2.99, 4, 8.54, 13.17, 17.85, 22.43, 26.99, 31.57, 36.14, 
    40.82, 45.44, 50.02 ;

 PG1 = 0.09, 0.88, 1.86, 2.84, 7.49, 12.05, 16.61, 21.28, 25.9, 30.43, 35.03, 
    39.65, 44.33, 48.84 ;

 PG15 = 0.06, 0.86, 1.87, 2.84, 7.48, 12.03, 16.65, 21.29, 25.86, 30.46, 
    35.02, 39.66, 44.3, 48.9 ;

 PG30 = 0.09, 0.85, 1.86, 2.85, 7.49, 12.01, 16.66, 21.31, 25.87, 30.43, 
    35.05, 39.71, 44.32, 48.87 ;

 PG60 = 0.09, 0.85, 1.85, 2.84, 7.49, 12.04, 16.68, 21.31, 25.87, 30.43, 
    35.05, 39.7, 44.31, 48.83 ;

 V1 = 23, 48, 121, 125, 130, 132, 133, 133, 133, 135, 135, 135, 135, 137 ;

 V15 = 32, 72, 123, 126, 130, 132, 133, 133, 133, 135, 135, 135, 135, 136 ;

 V30 = 36, 89, 123, 126, 130, 132, 133, 134, 134, 134, 135, 135, 136, 136 ;

 V60 = 39, 111, 123, 126, 130, 132, 133, 133, 134, 134, 135, 135, 135, 135 ;

 CREEP = 3, 22, 0, 0, 0, 0, 0, -1, 0, 0, 0, 0, -1, -1 ;

 DELT60 = 39, 72, 12, 3, 4, 2, 1, 0, 1, 0, 1, 0, 0, 0 ;
}
