netcdf data {
dimensions:
	time = UNLIMITED ; // (976 currently)
variables:
	float time(time) ;
		time:unit = "s" ;
		time:label = "Temps" ;
	float DEPTH(time) ;
		DEPTH:unit = "m" ;
		DEPTH:label = "Prof." ;
	float AS(time) ;
		AS:unit = "m/h" ;
		AS:label = "VIA" ;
		AS:scale_max = 1500.f ;
	int EVP(time) ;
		EVP:label = "evt-part" ;
	int EVR(time) ;
		EVR:label = "evt-new-rod" ;
	float TP(time) ;
		TP:unit = "bar" ;
		TP:label = "PO" ;
		TP:scale_max = 300.f ;
	float IP(time) ;
		IP:unit = "bar" ;
		IP:label = "PI" ;
		IP:scale_max = 50.f ;
	float TQ(time) ;
		TQ:unit = "bar" ;
		TQ:label = "CR" ;
		TQ:scale_max = 300.f ;
	float SP(time) ;
		SP:unit = "bar" ;
		SP:label = "PF" ;
		SP:scale_max = 300.f ;
data:

 time = 0, 2.2, 2.4, 2.6, 2.8, 3, 3.2, 3.4, 3.6, 3.8, 4, 4.2, 4.4, 4.6, 4.8, 
    5, 5.2, 5.4, 5.6, 5.8, 29, 29.2, 29.4, 29.6, 29.8, 30.2, 30.6, 31.2, 
    31.8, 32.8, 33.6, 34.4, 35.6, 36.8, 37.6, 38.2, 38.8, 39.4, 39.8, 40.2, 
    40.4, 40.6, 40.8, 41, 41.2, 41.4, 41.6, 41.8, 42.2, 42.6, 42.8, 89.2, 
    89.6, 90.2, 91.2, 93.4, 94.2, 115.8, 118.2, 119, 119.8, 120.4, 122.4, 
    125.6, 128.2, 130.399, 131, 131.4, 131.8, 132.2, 132.4, 132.6, 133, 
    133.4, 133.8, 134.2, 134.4, 134.8, 135, 135.2, 135.4, 135.6, 135.8, 136, 
    136.2, 136.4, 136.6, 136.8, 137.2, 137.8, 148.2, 158.6, 165.8, 173.6, 
    178.8, 183.4, 192.8, 197.2, 205.6, 215.4, 221.6, 228.6, 236, 245.2, 252, 
    256.799, 263, 269.6, 276.8, 284, 289.6, 297, 303.8, 308.8, 317.4, 323.8, 
    329.8, 331.6, 334, 338.2, 341.8, 345, 347.2, 349.8, 351, 352.8, 354, 
    354.4, 354.6, 354.8, 355, 355.2, 355.4, 355.6, 355.8, 356, 356.2, 356.4, 
    356.6, 356.8, 357, 357.2, 357.4, 357.6, 359.8, 360, 425.2, 425.4, 425.6, 
    426, 427, 428.2, 430.2, 432.2, 434.8, 436, 438.8, 439.8, 441, 443, 444.8, 
    445.8, 448.6, 451.8, 454.2, 458.8, 462.2, 464.2, 465.4, 466.2, 467.8, 
    468.6, 469.6, 470.2, 470.8, 471.4, 472, 473.2, 474, 474.6, 475.2, 475.8, 
    476.6, 477.2, 478, 478.6, 479, 479.4, 480.2, 480.6, 481.4, 482.6, 483.4, 
    484.2, 484.6, 485.2, 485.6, 487, 488, 489.4, 490.6, 492.8, 496.2, 498.2, 
    500.6, 504.4, 506.8, 508.8, 510.8, 513.599, 515.8, 517.8, 519.4, 521.4, 
    524, 527, 528.6, 529.8, 530.8, 531.6, 534.2, 535.4, 536.8, 538, 539.2, 
    539.8, 541.2, 543, 557.4, 587.8, 608.2, 640.8, 661.2, 674.6, 1066.8, 
    1096.4, 1121, 1144, 1168.4, 1178.6, 1184.6, 1188.4, 1190, 1191.2, 1191.8, 
    1192.4, 1193, 1194.2, 1195.4, 1197.8, 1204.2, 1206.4, 1207.4, 1209, 
    1210.8, 1212.4, 1213.8, 1214.8, 1215.4, 1216, 1216.8, 1217.8, 1219.6, 
    1220.6, 1221.8, 1222.6, 1223.6, 1224.2, 1225, 1225.8, 1227.4, 1228.6, 
    1230, 1231, 1231.8, 1232.4, 1233.6, 1234.2, 1235.8, 1236.4, 1237, 1238.8, 
    1240.6, 1243, 1247.4, 1249, 1251.4, 1254.2, 1258.4, 1263.4, 1268.6, 
    1272.8, 1275.4, 1277, 1278.6, 1279.2, 1279.8, 1280.4, 1281.2, 1290, 
    1291.4, 1293, 1293.6, 1294.2, 1294.6, 1296.4, 1303.6, 1306.8, 1308.4, 
    1310.4, 1312.4, 1314, 1359.6, 1360.6, 1362, 1362.6, 1363.2, 1363.8, 
    1364.4, 1365, 1365.4, 1366, 1366.8, 1367.4, 1368, 1368.8, 1369.6, 1370.4, 
    1372, 1373.6, 1375, 1376.8, 1377.6, 1378.2, 1378.6, 1379, 1379.4, 1379.6, 
    1379.8, 1380, 1380.2, 1380.4, 1380.6, 1380.8, 1381, 1381.2, 1381.4, 
    1381.6, 1381.8, 1382, 1382.2, 1382.4, 1382.8, 1383.2, 1383.6, 1384, 
    1384.4, 1384.6, 1384.8, 1385, 1385.2, 1385.4, 1385.6, 1385.8, 1386, 
    1386.2, 1386.4, 1386.6, 1386.8, 1387, 1387.2, 1387.4, 1387.6, 1387.8, 
    1388, 1388.2, 1388.4, 1388.6, 1388.8, 1389.2, 1390.4, 1393, 1395, 1396.2, 
    1399.2, 1402.8, 1408, 1410.4, 1414.6, 1420, 1425.8, 1428.6, 1431.8, 
    1437.6, 1443, 1450.4, 1452.8, 1457.6, 1463.4, 1466, 1472.4, 1476.6, 1481, 
    1485.6, 1491.2, 1495, 1498, 1862.8, 1863.4, 1865, 1866.2, 1868.2, 1870, 
    1872.6, 1876.2, 1878.8, 1880.8, 1882.4, 1883.8, 1885.4, 1889.6, 1892.2, 
    1897.8, 1900.8, 1905.2, 1907.6, 1912.8, 1915.2, 1918, 1920.2, 1922.8, 
    1925.4, 1928.2, 1931.2, 1933, 1935.8, 1938, 1942.4, 1948.4, 1951.4, 
    1952.2, 1953.6, 1955.6, 1959.2, 1960.8, 1962.2, 1963, 1964, 1965.4, 
    1967.2, 1969.6, 1971.4, 1972.2, 1974.6, 1975.8, 1978.6, 1981, 1984.8, 
    1987.2, 1989.6, 1991.4, 1992.8, 1995.2, 1997, 1999, 2000.2, 2003.8, 
    2005.6, 2007.4, 2009.4, 2011.6, 2013.6, 2014.4, 2015.2, 2016.6, 2017.4, 
    2018.8, 2020.2, 2022, 2023, 2024.6, 2026.6, 2028.6, 2029.8, 2031, 2031.6, 
    2032.2, 2032.6, 2033, 2033.4, 2033.8, 2034.2, 2034.6, 2035, 2035.4, 
    2035.8, 2036.6, 2037.2, 2037.8, 2038.2, 2039, 2040, 2041, 2041.6, 2043, 
    2045, 2046.6, 2048, 2049.2, 2050.6, 2052.2, 2054.399, 2055, 2055.399, 
    2055.6, 2056, 2056.2, 2056.399, 2056.6, 2056.8, 2057, 2057.2, 2057.399, 
    2057.6, 2057.8, 2058, 2060.8, 2066.6, 2075.8, 2079.6, 2085.399, 2363.2, 
    2372.8, 2383.4, 2385.4, 2389.4, 2391.6, 2393.4, 2395, 2396.4, 2398, 
    2399.6, 2401, 2402, 2403.6, 2405.2, 2407, 2408.4, 2410.6, 2412.8, 2414, 
    2482.2, 2483.2, 2484, 2485, 2486, 2486.8, 2487.6, 2488.6, 2489.6, 2490.4, 
    2491.8, 2493.2, 2494.6, 2495.8, 2497.4, 2498.8, 2500.6, 2501.4, 2502.8, 
    2504.2, 2505.6, 2507.4, 2509.6, 2511.6, 2513.2, 2515.2, 2517, 2518.4, 
    2518.8, 2519.2, 2527.6, 2534.2, 2537.4, 2542.6, 2550.8, 2558.4, 2565.2, 
    2573.8, 2583.8, 2590.6, 2596.6, 2600.4, 2602, 2602.6, 2603.2, 2604.4, 
    2605.8, 2608, 2608.4, 2608.8, 2609, 2609.2, 2609.4, 2609.8, 2610.4, 
    2612.6, 2614.6, 2616, 2617.2, 2617.8, 2618.6, 2619.4, 2620.2, 2622.2, 
    2625.2, 2629, 2631.6, 2633, 2634, 2634.4, 2637.8, 2638.4, 2639.2, 2639.8, 
    2641, 2643, 2645.2, 2652.6, 2662.2, 2668.8, 2673, 2682.6, 2757.2, 2767, 
    2777.6, 2780, 2782.4, 2783, 2784.2, 2787, 2790.4, 2794.8, 2802.8, 2803.4, 
    2805.4, 2806.4, 2808, 2809.6, 2811.8, 2814.4, 2817, 2823.2, 2825.4, 
    2828.4, 2833.4, 2842.2, 2852.2, 2854, 2855, 2857.8, 2860.6, 2864.6, 
    2870.4, 2871, 2872, 2873.2, 2875, 2876.6, 2877.4, 2878.2, 2878.6, 2879, 
    2879.4, 2880.2, 2885, 2888.8, 2891.6, 2896, 2897.8, 2898.8, 2900, 2901.4, 
    2902.6, 2904.4, 2906.2, 2908.8, 2910.4, 2916.2, 2919.8, 2920.4, 2921.4, 
    2923, 2923.6, 2924.8, 2926.2, 2926.8, 2928, 2929.2, 2930.2, 2931.4, 
    2932.8, 2933.4, 2934.2, 2935.8, 2937.6, 2941, 2941.6, 2941.8, 2942.4, 
    2943.2, 2944.8, 2948.6, 3063.4, 3064.8, 3066.6, 3068.6, 3071, 3073.8, 
    3076.8, 3087, 3090.8, 3094.2, 3095.6, 3096.2, 3097.2, 3098.8, 3100.2, 
    3101.8, 3103, 3104.6, 3107, 3112, 3114.2, 3116.8, 3117.8, 3118.6, 3119.2, 
    3120, 3120.4, 3121.8, 3122.8, 3126, 3127.6, 3129, 3131.2, 3133.8, 3137.8, 
    3139.4, 3140.8, 3141.8, 3142.8, 3143.8, 3145.4, 3146.8, 3148.2, 3149.2, 
    3150.4, 3151.4, 3152.8, 3155.2, 3157.6, 3158.8, 3159.8, 3161, 3162, 
    3163.2, 3163.8, 3164.2, 3165.8, 3174.2, 3176.8, 3177.6, 3178, 3179.8, 
    3186.2, 3190.4, 3194, 3199.6, 3203.6, 3210.8, 3215.2, 3220.8, 3228.2, 
    3235, 3241.2, 3247.6, 3251.2, 3253, 3259, 3266.2, 3272.4, 3277.8, 3592.8, 
    3595, 3596.4, 3597.4, 3599, 3600.8, 3605.2, 3609, 3610.4, 3612, 3613.4, 
    3614.6, 3618.2, 3619.4, 3620.6, 3621.8, 3624.4, 3625.8, 3627.4, 3630.4, 
    3631.8, 3633.4, 3634.8, 3636.2, 3638, 3639.6, 3641.2, 3643.8, 3645.6, 
    3647.4, 3649.4, 3651.4, 3653.2, 3655.4, 3656.8, 3657.2, 3657.4, 3657.8, 
    3680.4, 3683.4, 3688, 3693.4, 3698, 3704, 3708.2, 3712.4, 3714.4, 3718, 
    3721, 3724.6, 3727.4, 3730.2, 3733, 3736, 3741.6, 3746.2, 3752.2, 3755.8, 
    3762.2, 3765.6, 3767.8, 3769.4, 3769.8, 3770, 3770.4, 3770.8, 3774, 3783, 
    3787, 3789.6, 3791.4, 3792.6, 3793.8, 3795, 3796.2, 3798.4, 3799.8, 
    3800.4, 3801.2, 3801.8, 3802.8, 3805.4, 3854, 3855.2, 3857, 3858.6, 
    3860.8, 3863.4, 3866, 3867.2, 3869.6, 3870.4, 3871.6, 3873.2, 3874.8, 
    3880.8, 3891.8, 3900.2, 3908.6, 3917.8, 3926, 3930.4, 3932, 3932.6, 
    3933.2, 3934, 3934.6, 3935.2, 3935.8, 3936.4, 3937.4, 3943.2, 3946, 
    3946.4, 3946.8, 3947.4, 3949, 3951.6, 3952, 3952.4, 3953.8, 3954.2, 
    3954.6, 3955.2, 3956.2, 3956.6, 3957, 3957.2, 3957.6, 3958.2, 3958.8, 
    3959.2, 3959.6, 3960, 3963.6, 3964.2, 3965, 3966.2, 3966.8, 3967.8, 3970, 
    3972.4, 3974.8, 3978, 3979.2, 3980.2, 3982.2, 3983.4, 3984, 3985.8, 
    3986.8, 3988.4, 3991.4, 3992.2, 3993.6, 3994.8, 3995.6, 3998.4, 3999.8, 
    4001.2, 4002.8, 4004.4, 4005.8, 4007.4, 4009, 4010.4, 4012.2, 4013.4, 
    4015.4, 4017.6, 4019, 4020.6, 4022.8, 4024, 4027.2, 4028.8, 4032.8, 
    4037.6, 4042.4, 4043.6, 4046, 4047, 4163.4 ;

 DEPTH = 0, 0.02, 0.08, 0.15, 0.21, 0.28, 0.35, 0.42, 0.48, 0.55, 0.62, 0.69, 
    0.76, 0.83, 0.9, 0.97, 1.04, 1.11, 1.19, 1.24, 1.25, 1.27, 1.28, 1.29, 
    1.3, 1.32, 1.33, 1.34, 1.35, 1.37, 1.38, 1.39, 1.4, 1.41, 1.42, 1.44, 
    1.45, 1.46, 1.47, 1.5, 1.52, 1.53, 1.54, 1.56, 1.57, 1.59, 1.6, 1.61, 
    1.63, 1.65, 1.66, 1.67, 1.69, 1.7, 1.71, 1.72, 1.73, 1.75, 1.76, 1.77, 
    1.78, 1.79, 1.8, 1.81, 1.82, 1.83, 1.85, 1.86, 1.87, 1.89, 1.9, 1.91, 
    1.92, 1.94, 1.95, 1.97, 1.98, 2, 2.01, 2.03, 2.05, 2.07, 2.08, 2.09, 
    2.11, 2.12, 2.13, 2.14, 2.16, 2.17, 2.19, 2.2, 2.21, 2.22, 2.23, 2.24, 
    2.26, 2.27, 2.28, 2.29, 2.31, 2.32, 2.33, 2.34, 2.35, 2.36, 2.37, 2.38, 
    2.4, 2.41, 2.42, 2.43, 2.45, 2.46, 2.47, 2.48, 2.49, 2.5, 2.51, 2.53, 
    2.54, 2.55, 2.56, 2.57, 2.58, 2.59, 2.61, 2.62, 2.65, 2.69, 2.75, 2.81, 
    2.88, 2.95, 3.02, 3.09, 3.16, 3.23, 3.3, 3.36, 3.43, 3.5, 3.56, 3.61, 
    3.64, 3.66, 3.68, 3.7, 3.71, 3.73, 3.74, 3.75, 3.77, 3.78, 3.79, 3.8, 
    3.82, 3.83, 3.84, 3.85, 3.87, 3.88, 3.89, 3.91, 3.92, 3.93, 3.95, 3.96, 
    3.97, 3.98, 3.99, 4, 4.01, 4.02, 4.04, 4.05, 4.06, 4.07, 4.08, 4.1, 4.11, 
    4.12, 4.13, 4.15, 4.16, 4.17, 4.19, 4.2, 4.21, 4.22, 4.24, 4.25, 4.26, 
    4.27, 4.28, 4.3, 4.31, 4.33, 4.34, 4.35, 4.36, 4.37, 4.39, 4.4, 4.41, 
    4.43, 4.44, 4.45, 4.46, 4.47, 4.49, 4.5, 4.51, 4.53, 4.54, 4.55, 4.57, 
    4.58, 4.6, 4.61, 4.62, 4.63, 4.64, 4.65, 4.66, 4.67, 4.68, 4.69, 4.7, 
    4.71, 4.72, 4.74, 4.75, 4.76, 4.77, 4.78, 4.79, 4.8, 4.82, 4.83, 4.84, 
    4.85, 4.86, 4.87, 4.89, 4.91, 4.92, 4.93, 4.94, 4.95, 4.97, 4.98, 5, 
    5.01, 5.02, 5.03, 5.05, 5.06, 5.08, 5.09, 5.1, 5.11, 5.12, 5.13, 5.15, 
    5.16, 5.18, 5.19, 5.2, 5.21, 5.24, 5.25, 5.26, 5.27, 5.28, 5.29, 5.31, 
    5.32, 5.33, 5.34, 5.36, 5.37, 5.38, 5.39, 5.4, 5.41, 5.43, 5.44, 5.45, 
    5.47, 5.48, 5.49, 5.5, 5.51, 5.52, 5.53, 5.54, 5.56, 5.57, 5.58, 5.6, 
    5.61, 5.62, 5.64, 5.65, 5.66, 5.67, 5.68, 5.69, 5.71, 5.72, 5.73, 5.74, 
    5.75, 5.77, 5.78, 5.79, 5.81, 5.82, 5.83, 5.84, 5.85, 5.87, 5.88, 5.89, 
    5.9, 5.92, 5.93, 5.94, 5.95, 5.96, 5.98, 5.99, 6, 6.02, 6.04, 6.06, 6.07, 
    6.08, 6.1, 6.11, 6.13, 6.14, 6.16, 6.18, 6.2, 6.22, 6.24, 6.26, 6.28, 
    6.29, 6.3, 6.32, 6.33, 6.34, 6.36, 6.38, 6.4, 6.44, 6.47, 6.5, 6.53, 
    6.55, 6.59, 6.64, 6.69, 6.74, 6.8, 6.85, 6.91, 6.97, 7.02, 7.07, 7.13, 
    7.19, 7.25, 7.3, 7.33, 7.34, 7.36, 7.38, 7.39, 7.41, 7.42, 7.43, 7.45, 
    7.47, 7.48, 7.49, 7.51, 7.52, 7.53, 7.54, 7.56, 7.57, 7.58, 7.59, 7.61, 
    7.62, 7.63, 7.64, 7.66, 7.67, 7.68, 7.7, 7.71, 7.73, 7.74, 7.75, 7.77, 
    7.78, 7.79, 7.8, 7.81, 7.83, 7.84, 7.85, 7.86, 7.87, 7.88, 7.9, 7.91, 
    7.92, 7.93, 7.95, 7.96, 7.98, 7.99, 8.01, 8.02, 8.03, 8.05, 8.06, 8.08, 
    8.09, 8.11, 8.12, 8.13, 8.14, 8.15, 8.16, 8.18, 8.19, 8.2, 8.21, 8.23, 
    8.24, 8.25, 8.26, 8.28, 8.29, 8.3, 8.31, 8.33, 8.34, 8.35, 8.37, 8.38, 
    8.4, 8.41, 8.43, 8.44, 8.45, 8.47, 8.48, 8.49, 8.51, 8.52, 8.54, 8.55, 
    8.56, 8.58, 8.59, 8.6, 8.61, 8.62, 8.64, 8.65, 8.66, 8.67, 8.68, 8.7, 
    8.71, 8.73, 8.74, 8.76, 8.77, 8.78, 8.8, 8.82, 8.83, 8.84, 8.86, 8.87, 
    8.89, 8.9, 8.92, 8.93, 8.94, 8.96, 8.97, 8.98, 8.99, 9, 9.02, 9.03, 9.05, 
    9.06, 9.07, 9.08, 9.09, 9.11, 9.12, 9.14, 9.15, 9.17, 9.18, 9.2, 9.22, 
    9.24, 9.26, 9.29, 9.31, 9.35, 9.38, 9.4, 9.42, 9.43, 9.44, 9.45, 9.46, 
    9.47, 9.48, 9.49, 9.5, 9.51, 9.52, 9.54, 9.55, 9.56, 9.57, 9.58, 9.6, 
    9.61, 9.62, 9.63, 9.65, 9.66, 9.67, 9.69, 9.7, 9.71, 9.72, 9.73, 9.75, 
    9.76, 9.77, 9.78, 9.8, 9.81, 9.82, 9.83, 9.84, 9.85, 9.86, 9.88, 9.89, 
    9.9, 9.91, 9.92, 9.93, 9.94, 9.95, 9.97, 9.98, 9.99, 10, 10.01, 10.02, 
    10.03, 10.05, 10.06, 10.07, 10.08, 10.09, 10.1, 10.11, 10.12, 10.14, 
    10.15, 10.16, 10.18, 10.19, 10.2, 10.21, 10.22, 10.23, 10.24, 10.26, 
    10.27, 10.28, 10.29, 10.31, 10.32, 10.33, 10.34, 10.36, 10.37, 10.38, 
    10.39, 10.4, 10.41, 10.43, 10.44, 10.45, 10.46, 10.47, 10.48, 10.5, 
    10.51, 10.52, 10.53, 10.54, 10.55, 10.56, 10.58, 10.59, 10.6, 10.61, 
    10.63, 10.64, 10.65, 10.66, 10.67, 10.68, 10.69, 10.7, 10.72, 10.73, 
    10.74, 10.75, 10.76, 10.77, 10.79, 10.8, 10.82, 10.83, 10.84, 10.85, 
    10.86, 10.87, 10.89, 10.9, 10.91, 10.92, 10.94, 10.95, 10.96, 10.97, 
    10.98, 11, 11.01, 11.03, 11.04, 11.05, 11.06, 11.08, 11.09, 11.1, 11.11, 
    11.12, 11.14, 11.15, 11.16, 11.17, 11.19, 11.2, 11.21, 11.23, 11.24, 
    11.25, 11.26, 11.27, 11.29, 11.3, 11.31, 11.32, 11.33, 11.34, 11.36, 
    11.37, 11.38, 11.39, 11.4, 11.42, 11.43, 11.45, 11.46, 11.47, 11.49, 
    11.51, 11.52, 11.53, 11.54, 11.56, 11.57, 11.59, 11.6, 11.61, 11.62, 
    11.64, 11.65, 11.67, 11.68, 11.69, 11.7, 11.71, 11.73, 11.74, 11.75, 
    11.76, 11.77, 11.79, 11.8, 11.81, 11.82, 11.84, 11.85, 11.86, 11.87, 
    11.88, 11.89, 11.91, 11.92, 11.94, 11.95, 11.96, 11.98, 11.99, 12, 12.01, 
    12.02, 12.03, 12.04, 12.06, 12.07, 12.08, 12.09, 12.1, 12.12, 12.13, 
    12.14, 12.15, 12.16, 12.18, 12.19, 12.2, 12.21, 12.23, 12.24, 12.25, 
    12.26, 12.27, 12.29, 12.3, 12.31, 12.33, 12.34, 12.35, 12.36, 12.38, 
    12.39, 12.4, 12.41, 12.42, 12.43, 12.45, 12.46, 12.47, 12.48, 12.49, 
    12.5, 12.51, 12.53, 12.54, 12.55, 12.56, 12.57, 12.58, 12.59, 12.61, 
    12.62, 12.64, 12.65, 12.67, 12.68, 12.69, 12.7, 12.71, 12.72, 12.73, 
    12.75, 12.76, 12.77, 12.78, 12.8, 12.82, 12.83, 12.84, 12.86, 12.87, 
    12.88, 12.9, 12.91, 12.92, 12.94, 12.95, 12.96, 12.98, 12.99, 13, 13.02, 
    13.03, 13.04, 13.05, 13.07, 13.08, 13.09, 13.11, 13.12, 13.13, 13.14, 
    13.16, 13.17, 13.18, 13.19, 13.21, 13.22, 13.23, 13.24, 13.25, 13.27, 
    13.28, 13.29, 13.3, 13.31, 13.32, 13.33, 13.34, 13.35, 13.37, 13.38, 
    13.39, 13.4, 13.41, 13.43, 13.44, 13.46, 13.47, 13.48, 13.49, 13.5, 
    13.51, 13.52, 13.53, 13.55, 13.56, 13.58, 13.59, 13.6, 13.62, 13.63, 
    13.64, 13.66, 13.67, 13.68, 13.7, 13.71, 13.72, 13.73, 13.75, 13.76, 
    13.78, 13.79, 13.8, 13.81, 13.82, 13.83, 13.85, 13.86, 13.87, 13.88, 
    13.89, 13.9, 13.92, 13.93, 13.94, 13.95, 13.97, 13.98, 13.99, 14.01, 
    14.02, 14.04, 14.05, 14.06, 14.08, 14.09, 14.11, 14.12, 14.14, 14.15, 
    14.17, 14.18, 14.19, 14.2, 14.22, 14.23, 14.24, 14.26, 14.27, 14.29, 
    14.3, 14.32, 14.33, 14.35, 14.36, 14.38, 14.39, 14.4, 14.42, 14.43, 
    14.44, 14.46, 14.47, 14.48, 14.49, 14.5, 14.51, 14.53, 14.54, 14.55, 
    14.57, 14.58, 14.59, 14.61, 14.62, 14.63, 14.64, 14.65, 14.67, 14.69, 
    14.7, 14.72, 14.73, 14.74, 14.76, 14.77, 14.78, 14.8, 14.81, 14.82, 
    14.84, 14.85, 14.86, 14.87, 14.88, 14.9, 14.91, 14.92, 14.93, 14.94, 
    14.96, 14.97, 14.98, 15 ;

 AS = 0, 31.45398, 1178.385, 1148.298, 1138.269, 1228.529, 1258.615, 
    1208.471, 1193.428, 1228.529, 1278.673, 1228.529, 1193.428, 1273.658, 
    1328.817, 1268.644, 1238.557, 1288.701, 1333.831, 882.5349, 1.642649, 
    340.9794, 320.9218, 180.5185, 195.5617, 135.3889, 110.3169, 68.53017, 
    70.20164, 40.11522, 47.63682, 46.38322, 40.95095, 35.93655, 48.89042, 
    83.57337, 75.21603, 78.55898, 92.76645, 220.6337, 330.9506, 240.6913, 
    240.6913, 260.7489, 245.7057, 265.7633, 240.6913, 220.6337, 180.5185, 
    155.4465, 185.5329, 1.210373, 97.78085, 70.20164, 39.11234, 25.07201, 
    48.89042, 2.367912, 15.04321, 48.89042, 46.38322, 60.17283, 19.55617, 
    13.47621, 14.65748, 18.23419, 85.24484, 100.288, 125.3601, 167.9825, 
    185.5329, 190.5473, 107.8097, 100.288, 125.3601, 167.9825, 180.5185, 
    205.5905, 215.6193, 325.9362, 335.965, 310.8929, 230.6625, 225.6481, 
    255.7345, 280.8065, 215.6193, 180.5185, 127.8673, 75.21603, 4.821541, 
    3.760802, 7.243026, 5.271551, 8.100188, 8.284665, 5.121092, 8.433313, 
    4.41745, 5.321407, 7.278971, 5.157671, 6.776219, 5.450438, 5.751815, 
    7.730537, 5.984932, 5.622209, 7.382315, 5.710847, 6.805261, 4.878878, 
    7.226639, 7.220739, 4.781175, 6.111303, 7.521604, 20.05761, 16.29681, 
    12.6554, 10.86454, 11.28241, 25.52787, 15.42893, 30.08641, 22.28623, 
    45.96535, 115.3313, 461.325, 722.074, 1027.953, 1198.442, 1303.745, 
    1218.5, 1193.428, 1238.557, 1268.644, 1253.601, 1213.485, 1218.5, 
    1278.673, 1208.471, 1123.226, 857.4628, 48.77646, 421.2098, 1.015186, 
    285.821, 200.5761, 152.9393, 45.12962, 46.80109, 27.07777, 21.06049, 
    17.35755, 31.75788, 19.69944, 36.1037, 35.93655, 22.56481, 25.62917, 
    39.11234, 20.05761, 16.29681, 19.63974, 10.24682, 15.33817, 22.06337, 
    31.75788, 47.63682, 23.81841, 45.12962, 42.12098, 61.8443, 61.8443, 
    70.20164, 60.17283, 32.59362, 73.96243, 71.8731, 76.8875, 65.18723, 
    57.66563, 75.21603, 65.18723, 90.25925, 110.3169, 127.8673, 45.12962, 
    110.3169, 58.91923, 42.62242, 45.12962, 50.14402, 102.7952, 75.21603, 
    135.3889, 40.11522, 42.12098, 32.23544, 36.77229, 18.69005, 13.56838, 
    20.05761, 19.22188, 16.09887, 15.04321, 18.05185, 20.55905, 19.34127, 
    18.23419, 26.07489, 30.71321, 22.56481, 17.35755, 17.71756, 32.59362, 
    47.63682, 45.12962, 55.15843, 14.65748, 32.59362, 25.78835, 30.92215, 
    30.92215, 63.51577, 28.65373, 21.17192, 2.64649, 1.187622, 1.868111, 
    1.261291, 1.81895, 2.694306, 1.439771, 1.21972, 1.46763, 1.61333, 
    1.97288, 4.031186, 7.18731, 10.29272, 23.81841, 38.44375, 101.9595, 
    105.3025, 83.57337, 31.75788, 32.59362, 15.46107, 8.148404, 25.98372, 
    43.12386, 23.81841, 26.18632, 30.71321, 32.23544, 56.16131, 81.90191, 
    65.18723, 52.65123, 39.11234, 27.30064, 40.11522, 41.78669, 62.68003, 
    53.15267, 70.20164, 50.14402, 68.94804, 48.89042, 30.08641, 40.11522, 
    36.1037, 46.38322, 60.17283, 42.62242, 63.51577, 22.56481, 90.25925, 
    91.93071, 22.28623, 25.07201, 15.87894, 10.0288, 23.19161, 17.13254, 
    14.32686, 11.93905, 10.63053, 7.328742, 8.596119, 18.12899, 26.32561, 
    23.19161, 76.8875, 63.51577, 65.18723, 68.94804, 4.786475, 39.39888, 
    25.69881, 63.51577, 95.27364, 95.27364, 20.61477, 6.825159, 12.84941, 
    26.95241, 21.56193, 24.57057, 24.44521, 0.9676917, 38.10946, 33.66813, 
    68.53017, 76.8875, 88.58778, 66.8587, 85.24484, 100.288, 71.8731, 
    67.69444, 78.55898, 61.8443, 56.41203, 53.90483, 47.63682, 30.08641, 
    23.81841, 31.5191, 28.9721, 53.90483, 81.90191, 122.8529, 175.5041, 
    193.0545, 235.6769, 245.7057, 215.6193, 290.8354, 245.7057, 270.7777, 
    325.9362, 366.0514, 366.0514, 356.0226, 376.0802, 406.1666, 300.8641, 
    230.6625, 195.5617, 122.8529, 112.8241, 132.8817, 92.76645, 190.5473, 
    486.397, 586.6851, 666.9155, 571.6419, 406.1666, 461.325, 686.9731, 
    827.3764, 972.7941, 957.7509, 972.7941, 972.7941, 1017.924, 1027.953, 
    962.7653, 972.7941, 1042.996, 1088.125, 1037.981, 867.4916, 556.5987, 
    265.7633, 130.3745, 52.65123, 18.51472, 31.08929, 39.27949, 18.72044, 
    16.71467, 12.53601, 15.46107, 11.22271, 9.471649, 6.397686, 15.04321, 
    11.90921, 10.20172, 7.614463, 5.014402, 19.22188, 10.86454, 7.089328, 
    16.97182, 7.678304, 13.37174, 9.345023, 10.90088, 11.10332, 11.6123, 
    17.04897, 0.1209615, 86.91631, 26.95241, 33.42935, 18.05185, 25.62917, 
    17.35755, 12.81458, 13.88604, 22.56481, 27.57921, 26.5047, 23.81841, 
    12.17783, 16.5861, 9.491548, 13.03745, 11.39637, 19.63974, 10.60739, 
    18.38614, 22.92298, 23.24859, 18.12899, 20.82906, 21.13212, 21.39478, 
    25.07201, 13.96869, 17.32248, 12.08015, 6.518723, 13.70603, 46.38322, 
    30.80276, 18.05185, 13.9289, 33.84722, 27.22104, 52.65123, 38.10946, 
    33.66813, 35.10082, 19.22188, 25.07201, 50.14402, 18.38614, 35.10082, 
    17.55041, 21.31121, 14.25146, 23.81841, 23.81841, 25.62917, 29.37007, 
    25.07201, 30.08641, 19.55617, 37.60802, 16.15752, 29.52926, 26.18632, 
    19.55617, 28.263, 21.06049, 46.38322, 47.63682, 32.23544, 61.42643, 
    32.23544, 40.11522, 20.05761, 36.1037, 25.07201, 28.58209, 25.57345, 
    41.78669, 47.63682, 85.24484, 88.58778, 90.25925, 147.9249, 160.4609, 
    97.78085, 132.8817, 132.8817, 160.4609, 137.8961, 130.3745, 72.70884, 
    85.24484, 61.8443, 95.27364, 53.90483, 44.12674, 42.12098, 80.23044, 
    40.83156, 24.06913, 28.83282, 35.81716, 30.08641, 28.65373, 23.81841, 
    26.43958, 75.21603, 185.5329, 215.6193, 172.9969, 215.6193, 305.8785, 
    351.0082, 381.0946, 376.0802, 396.1378, 521.4979, 636.8291, 571.6419, 
    371.0658, 18.26675, 6.916417, 4.36035, 9.500973, 7.608059, 2.259236, 
    4.178668, 3.406009, 18.55329, 9.527365, 17.32248, 22.84339, 23.19161, 
    32.95179, 30.71321, 25.07201, 32.95179, 36.1037, 35.10082, 25.69881, 
    30.64357, 27.22104, 25.07201, 20.96932, 35.10082, 0.6029047, 39.11234, 
    60.17283, 46.1325, 55.15843, 45.12962, 45.12962, 46.1325, 42.12098, 
    48.89042, 32.95179, 31.5191, 26.5047, 33.42935, 30.08641, 32.23544, 
    20.05761, 45.12962, 25.78835, 30.08641, 30.08641, 20.05761, 23.24859, 
    18.55329, 22.56481, 18.55329, 20.61477, 34.38448, 97.78085, 125.3601, 
    5.253183, 5.77416, 12.22261, 6.943019, 4.647495, 5.014402, 6.04678, 
    5.8307, 4.914114, 6.784192, 7.18731, 13.1958, 26.32561, 61.8443, 
    70.20164, 30.08641, 27.93739, 18.23419, 92.76645, 137.8961, 215.6193, 
    220.6337, 210.6049, 120.3457, 71.8731, 22.79274, 20.05761, 27.93739, 
    32.59362, 66.8587, 56.41203, 58.91923, 45.12962, 20.05761, 13.37174, 
    12.66796, 16.97182, 35.81716, 37.10658, 100.288, 11.20866, 60.17283, 
    48.89042, 65.18723, 40.95095, 27.57921, 16.41077, 5.014402, 5.536736, 
    6.230015, 8.596119, 3.969735, 0.4839638, 4.912068, 3.500621, 16.71467, 
    19.22188, 70.20164, 35.10082, 15.40138, 11.79859, 8.889168, 7.145524, 
    75.21603, 30.58785, 47.13538, 23.19161, 25.07201, 17.32248, 14.27176, 
    19.67189, 7.764236, 17.77834, 14.04033, 8.424196, 4.558547, 4.914114, 
    23.40055, 38.10946, 22.20664, 15.04321, 14.04033, 8.645521, 61.8443, 
    44.12674, 38.44375, 22.28623, 22.56481, 47.63682, 52.65123, 137.8961, 
    132.8817, 95.27364, 56.41203, 11.07347, 10.29272, 15.75955, 11.85222, 
    26.18632, 45.12962, 39.27949, 25.78835, 35.10082, 26.74348, 21.17192, 
    13.88604, 25.69881, 8.12679, 10.30738, 68.53017, 47.13538, 27.57921, 
    70.20164, 35.10082, 49.42768, 70.20164, 46.80109, 38.44375, 58.16707, 
    45.12962, 33.66813, 70.20164, 62.68003, 30.08641, 26.74348, 15.9281, 
    70.20164, 200.5761, 75.21603, 61.42643, 36.35442, 14.51538, 0.3406998, 
    36.5335, 20.05761, 19.05473, 20.89334, 14.32686, 16.04609, 3.6379, 
    11.6123, 13.27342, 33.66813, 65.18723, 48.13826, 29.45961, 35.10082, 
    26.32561, 35.93655, 23.19161, 15.87894, 13.4386, 17.32248, 18.51472, 
    40.11522, 62.68003, 75.21603, 55.15843, 90.25925, 29.37007, 36.1037, 
    15.04321, 28.83282, 31.5191, 23.24859, 16.5861, 9.025925, 23.19161, 
    29.37007, 42.12098, 52.14978, 47.13538, 23.81841, 30.80276, 28.65373, 
    40.11522, 40.11522, 49.14114, 30.80276, 16.71467, 18.38614, 32.59362, 
    45.12962, 34.26508, 48.13826, 51.81549, 88.58778, 90.25925, 25.07201, 
    6.088917, 15.04321, 48.89042, 100.288, 21.17192, 7.678304, 9.551243, 
    11.70027, 6.626175, 9.025925, 6.407292, 10.0288, 7.163432, 6.098598, 
    6.04678, 5.984932, 8.148404, 10.30738, 23.9577, 6.017283, 5.989425, 
    9.54354, 10.21452, 0.1814736, 18.69005, 28.65373, 37.10658, 24.44521, 
    26.18632, 8.205386, 12.14013, 29.37007, 35.72762, 27.93739, 37.60802, 
    15.32178, 45.12962, 41.78669, 40.95095, 22.75767, 31.5191, 26.32561, 
    14.70891, 30.08641, 32.59362, 40.11522, 31.5191, 22.28623, 32.59362, 
    28.20601, 20.44333, 25.62917, 21.72908, 27.57921, 22.56481, 24.51486, 
    20.05761, 27.22104, 165.4753, 195.5617, 112.8241, 1.86376, 16.38038, 
    11.33691, 7.800182, 8.284665, 8.691631, 10.26759, 9.790024, 18.05185, 
    13.37174, 13.70603, 10.58596, 14.68504, 15.04321, 13.25235, 12.36886, 
    8.237947, 7.84863, 7.18731, 11.14312, 5.797903, 13.56838, 17.77834, 
    29.45961, 130.3745, 195.5617, 150.4321, 92.76645, 12.84941, 4.79154, 
    10.78096, 14.65748, 25.07201, 32.59362, 41.78669, 37.60802, 49.30829, 
    25.07201, 30.08641, 81.90191, 50.14402, 76.8875, 46.1325, 24.68629, 
    0.7841452, 43.45816, 20.61477, 28.83282, 18.69005, 18.51472, 24.68629, 
    36.77229, 20.47548, 51.39762, 30.92215, 23.81841, 28.20601, 6.518723, 
    3.282154, 5.491965, 4.53684, 5.450438, 4.525192, 10.71259, 28.83282, 
    83.57337, 68.53017, 71.45524, 60.17283, 88.58778, 100.288, 65.18723, 
    46.1325, 9.164253, 16.11772, 147.9249, 137.8961, 71.8731, 32.59362, 
    21.21478, 152.9393, 120.3457, 37.24985, 90.25925, 110.3169, 108.6454, 
    43.12386, 100.288, 147.9249, 195.5617, 140.4033, 83.57337, 93.60218, 
    132.8817, 157.9537, 105.3025, 18.10756, 66.8587, 51.39762, 40.95095, 
    70.20164, 55.15843, 21.88103, 15.46107, 15.46107, 15.67001, 30.92215, 
    36.1037, 26.57633, 42.62242, 60.17283, 32.87219, 40.11522, 28.20601, 
    19.05473, 46.38322, 30.80276, 38.44375, 53.90483, 24.35567, 35.81716, 
    42.98059, 31.34002, 33.22042, 30.80276, 33.84722, 33.84722, 27.22104, 
    24.51486, 33.42935, 26.57633, 25.98372, 30.08641, 22.56481, 19.60176, 
    39.27949, 12.84941, 31.34002, 11.03169, 8.566271, 7.939471, 36.77229, 
    15.87894, 53.15267, 20.05761 ;

 EVP = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EVR = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TP = 7.42, 7.42, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 
    70.89, 70.89, 70.89, 70.89, 69.67, 69.67, 69.67, 67.23, 69.67, 69.67, 
    73.34, 70.89, 69.67, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 
    70.89, 72.12, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 
    70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 69.67, 70.89, 70.89, 
    70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 
    73.34, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 
    70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 
    70.89, 69.67, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 
    70.89, 70.89, 70.89, 70.89, 72.12, 70.89, 70.89, 72.12, 70.89, 70.89, 
    70.89, 73.34, 70.89, 72.12, 70.89, 73.34, 73.34, 70.89, 73.34, 73.34, 
    73.34, 73.34, 73.34, 70.89, 70.89, 70.89, 72.12, 73.34, 70.89, 70.89, 
    73.34, 73.34, 70.89, 73.34, 70.89, 73.34, 70.89, 70.89, 70.89, 67.23, 
    66.01, 64.79, 64.79, 56.25, 56.25, 56.25, 57.47, 53.8, 55.03, 55.03, 
    53.8, 63.57, 63.57, 66.01, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 
    73.34, 70.89, 70.89, 70.89, 70.89, 73.34, 70.89, 70.89, 69.67, 70.89, 
    69.67, 73.34, 70.89, 70.89, 70.89, 70.89, 70.89, 72.12, 73.34, 73.34, 
    70.89, 72.12, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 73.34, 
    73.34, 73.34, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 
    70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 
    73.34, 70.89, 70.89, 70.89, 73.34, 70.89, 73.34, 73.34, 70.89, 70.89, 
    70.89, 73.34, 73.34, 69.67, 70.89, 70.89, 70.89, 73.34, 73.34, 70.89, 
    70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 73.34, 73.34, 73.34, 
    72.12, 73.34, 73.34, 73.34, 70.89, 73.34, 70.89, 72.12, 70.89, 70.89, 
    70.89, 70.89, 73.34, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 
    61.13, 68.45, 70.89, 70.89, 70.89, 73.34, 73.34, 73.34, 72.12, 70.89, 
    72.12, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 
    70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 
    70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 
    73.34, 70.89, 70.89, 73.34, 69.67, 70.89, 69.67, 70.89, 70.89, 70.89, 
    70.89, 70.89, 69.67, 70.89, 70.89, 72.12, 70.89, 73.34, 70.89, 70.89, 
    72.12, 73.34, 73.34, 70.89, 70.89, 73.34, 70.89, 72.12, 70.89, 70.89, 
    70.89, 70.89, 70.89, 70.89, 72.12, 73.34, 73.34, 70.89, 70.89, 73.34, 
    70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 
    70.89, 70.89, 70.89, 70.89, 69.67, 70.89, 70.89, 69.67, 69.67, 70.89, 
    70.89, 70.89, 73.34, 72.12, 70.89, 70.89, 67.23, 67.23, 66.01, 66.01, 
    68.45, 70.89, 68.45, 67.23, 66.01, 66.01, 66.01, 66.01, 64.79, 66.01, 
    66.01, 66.01, 64.79, 64.79, 64.79, 66.01, 66.01, 68.45, 70.89, 70.89, 
    70.89, 70.89, 70.89, 70.89, 70.89, 73.34, 70.89, 70.89, 70.89, 70.89, 
    70.89, 70.89, 70.89, 70.89, 70.89, 73.34, 70.89, 70.89, 70.89, 70.89, 
    70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 
    70.89, 72.12, 73.34, 73.34, 70.89, 70.89, 73.34, 70.89, 73.34, 72.12, 
    70.89, 70.89, 73.34, 67.23, 70.89, 70.89, 70.89, 66.01, 70.89, 70.89, 
    70.89, 69.67, 70.89, 70.89, 70.89, 73.34, 70.89, 70.89, 70.89, 70.89, 
    70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 
    70.89, 70.89, 70.89, 72.12, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 
    70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 
    70.89, 70.89, 67.23, 70.89, 67.23, 70.89, 69.67, 69.67, 70.89, 72.12, 
    69.67, 70.89, 70.89, 70.89, 70.89, 69.67, 70.89, 70.89, 70.89, 70.89, 
    73.34, 70.89, 70.89, 70.89, 70.89, 70.89, 70.89, 69.67, 69.67, 72.12, 
    73.34, 70.89, 70.89, 70.89, 70.89, 73.34, 69.67, 73.34, 70.89, 70.89, 
    73.34, 70.89, 69.67, 70.89, 70.89, 70.89, 70.89, 70.89, 69.67, 69.67, 
    69.67, 70.89, 68.45, 66.01, 67.23, 70.89, 73.34, 73.34, 73.34, 70.89, 
    70.89, 73.34, 70.89, 73.34, 74.56, 72.12, 73.34, 73.34, 73.34, 73.34, 
    73.34, 73.34, 73.34, 73.34, 73.34, 73.34, 73.34, 73.34, 72.12, 73.34, 
    73.34, 70.89, 70.89, 73.34, 73.34, 73.34, 73.34, 70.89, 73.34, 73.34, 
    73.34, 73.34, 73.34, 73.34, 70.89, 72.12, 70.89, 73.34, 73.34, 73.34, 
    74.56, 73.34, 73.34, 74.56, 74.56, 70.89, 73.34, 73.34, 73.34, 73.34, 
    73.34, 72.12, 70.89, 73.34, 74.56, 73.34, 73.34, 70.89, 70.89, 73.34, 
    74.56, 73.34, 73.34, 73.34, 73.34, 73.34, 73.34, 70.89, 73.34, 70.89, 
    73.34, 70.89, 70.89, 70.89, 73.34, 73.34, 73.34, 70.89, 72.12, 73.34, 
    70.89, 70.89, 70.89, 73.34, 70.89, 73.34, 70.89, 73.34, 73.34, 73.34, 
    70.89, 73.34, 73.34, 70.89, 73.34, 73.34, 73.34, 70.89, 70.89, 73.34, 
    73.34, 73.34, 73.34, 73.34, 70.89, 73.34, 74.56, 73.34, 73.34, 70.89, 
    73.34, 73.34, 72.12, 73.34, 73.34, 70.89, 70.89, 73.34, 73.34, 73.34, 
    73.34, 73.34, 73.34, 70.89, 70.89, 73.34, 70.89, 72.12, 73.34, 73.34, 
    73.34, 72.12, 70.89, 70.89, 72.12, 73.34, 70.89, 73.34, 73.34, 70.89, 
    70.89, 70.89, 70.89, 70.89, 73.34, 69.67, 73.34, 73.34, 74.56, 74.56, 
    70.89, 73.34, 73.34, 73.34, 73.34, 70.89, 70.89, 73.34, 70.89, 70.89, 
    73.34, 73.34, 70.89, 70.89, 73.34, 70.89, 72.12, 73.34, 73.34, 73.34, 
    70.89, 70.89, 73.34, 73.34, 70.89, 74.56, 73.34, 73.34, 70.89, 73.34, 
    73.34, 73.34, 70.89, 74.56, 70.89, 74.56, 73.34, 74.56, 74.56, 73.34, 
    70.89, 73.34, 73.34, 73.34, 74.56, 70.89, 74.56, 73.34, 70.89, 74.56, 
    74.56, 74.56, 70.89, 70.89, 70.89, 73.34, 74.56, 73.34, 73.34, 73.34, 
    74.56, 70.89, 74.56, 74.56, 73.34, 73.34, 74.56, 74.56, 74.56, 73.34, 
    73.34, 74.56, 74.56, 73.34, 73.34, 74.56, 72.12, 74.56, 70.89, 73.34, 
    70.89, 73.34, 74.56, 74.56, 74.56, 73.34, 73.34, 73.34, 73.34, 72.12, 
    70.89, 74.56, 74.56, 70.89, 73.34, 73.34, 74.56, 73.34, 74.56, 73.34, 
    73.34, 74.56, 73.34, 73.34, 73.34, 73.34, 74.56, 74.56, 74.56, 74.56, 
    74.56, 73.34, 74.56, 74.56, 74.56, 73.34, 70.89, 73.34, 73.34, 73.34, 
    73.34, 73.34, 73.34, 72.12, 74.56, 63.57, 70.89, 74.56, 74.56, 70.89, 
    73.34, 73.34, 59.91, 74.56, 74.56, 74.56, 73.34, 74.56, 73.34, 73.34, 
    73.34, 74.56, 74.56, 73.34, 74.56, 73.34, 73.34, 74.56, 74.56, 74.56, 
    70.89, 74.56, 74.56, 73.34, 74.56, 74.56, 73.34, 73.34, 74.56, 73.34, 
    73.34, 74.56, 74.56, 73.34, 74.56, 74.56, 74.56, 73.34, 74.56, 73.34, 
    74.56, 74.56, 73.34, 74.56, 70.89, 74.56, 73.34, 74.56, 74.56, 74.56, 
    70.89, 73.34, 74.56, 73.34, 74.56, 74.56, 74.56, 73.34, 73.34, 73.34, 
    73.34, 74.56, 73.34, 74.56, 70.89, 70.89, 70.89, 74.56, 73.34, 73.34, 
    74.56, 72.12, 74.56, 73.34, 73.34, 74.56, 73.34, 74.56, 74.56, 74.56, 
    74.56, 73.34, 73.34, 74.56, 72.12, 70.89, 73.34, 74.56, 73.34, 73.34, 
    74.56, 73.34, 73.34, 74.56, 73.34, 74.56, 73.34, 74.56, 73.34, 73.34, 
    73.34, 74.56, 73.34, 73.34, 73.34, 74.56, 73.34, 73.34, 74.56, 74.56, 
    74.56, 73.34, 74.56, 73.34, 73.34, 73.34, 73.34, 72.12, 73.34, 74.56, 
    73.34, 73.34, 73.34, 74.56, 74.56, 74.56, 73.34, 74.56, 74.56, 74.56, 
    74.56, 73.34, 74.56, 73.34, 73.34, 70.89, 74.56, 73.34, 70.89, 74.56, 
    70.89, 73.34, 74.56, 74.56, 73.34, 73.34, 74.56, 74.56, 74.56, 74.56, 
    72.12, 73.34, 73.34, 74.56, 74.56, 73.34, 74.56, 72.12, 73.34, 74.56, 
    73.34, 74.56, 74.56, 74.56, 70.89, 4.98 ;

 IP = 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 
    1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 0.09, 1.31, 1.31, 0.09, 1.31, 1.31, 
    1.31, 1.31, 1.31, 0.09, 1.31, 1.31, 1.31, 1.31, 0.09, 1.31, 1.31, 0.09, 
    0.09, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 
    1.31, 0.09, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 17.18, 2.53, 1.31, 
    1.31, 1.31, 1.31, 0.09, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 0.09, 1.31, 
    1.31, 1.31, 1.31, 1.31, 1.31, 0.09, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 
    1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 4.98, 4.98, 2.53, 2.53, 1.31, 2.53, 
    1.31, 2.53, 1.31, 2.53, 1.31, 2.53, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 
    2.53, 1.31, 1.31, 1.31, 1.31, 2.53, 2.53, 1.31, 1.31, 2.53, 2.53, 1.31, 
    2.53, 1.31, 1.31, 1.31, 2.53, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 
    2.53, 1.31, 1.31, 1.31, 1.31, 1.31, 2.53, 1.31, 1.31, 1.31, 1.31, 1.31, 
    2.53, 2.53, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 2.53, 3.75, 
    7.42, 8.64, 17.18, 8.64, 4.98, 7.42, 7.42, 6.2, 7.42, 4.98, 14.74, 4.98, 
    4.98, 4.98, 7.42, 9.86, 17.18, 26.95, 8.64, 7.42, 12.3, 8.64, 4.98, 4.98, 
    7.42, 7.42, 8.64, 14.74, 20.84, 7.42, 4.98, 7.42, 8.64, 12.3, 20.84, 
    7.42, 12.3, 12.3, 8.64, 8.64, 12.3, 20.84, 17.18, 7.42, 7.42, 14.74, 
    11.08, 8.64, 7.42, 2.53, 2.53, 1.31, 2.53, 2.53, 1.31, 2.53, 3.75, 4.98, 
    12.3, 7.42, 7.42, 4.98, 4.98, 6.2, 18.4, 9.86, 7.42, 4.98, 4.98, 3.75, 
    2.53, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 
    1.31, 1.31, 1.31, 2.53, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 
    7.42, 6.2, 2.53, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 
    1.31, 2.53, 3.75, 4.98, 4.98, 6.2, 7.42, 12.3, 34.27, 31.83, 12.3, 12.3, 
    12.3, 7.42, 7.42, 7.42, 12.3, 6.2, 3.75, 6.2, 1.31, 1.31, 1.31, 1.31, 
    1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 
    1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 7.42, 1.31, 1.31, 1.31, 
    1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 
    1.31, 1.31, 2.53, 1.31, 2.53, 1.31, 2.53, 2.53, 2.53, 4.98, 6.2, 4.98, 
    2.53, 1.31, 1.31, 2.53, 2.53, 1.31, 1.31, 2.53, 1.31, 1.31, 1.31, 1.31, 
    1.31, 2.53, 2.53, 1.31, 1.31, 2.53, 1.31, 1.31, 1.31, 2.53, 1.31, 1.31, 
    1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 
    1.31, 2.53, 1.31, 1.31, 2.53, 1.31, 1.31, 1.31, 1.31, 1.31, 2.53, 2.53, 
    4.98, 7.42, 7.42, 2.53, 4.98, 4.98, 7.42, 4.98, 3.75, 8.64, 2.53, 7.42, 
    7.42, 6.2, 4.98, 4.98, 7.42, 6.2, 6.2, 7.42, 4.98, 7.42, 7.42, 7.42, 
    7.42, 1.31, 1.31, 1.31, 1.31, 2.53, 2.53, 7.42, 4.98, 4.98, 7.42, 4.98, 
    2.53, 2.53, 2.53, 1.31, 2.53, 2.53, 4.98, 7.42, 1.31, 2.53, 2.53, 3.75, 
    7.42, 12.3, 2.53, 4.98, 7.42, 3.75, 2.53, 4.98, 4.98, 2.53, 2.53, 2.53, 
    4.98, 7.42, 2.53, 2.53, 2.53, 2.53, 3.75, 3.75, 7.42, 2.53, 2.53, 2.53, 
    2.53, 2.53, 4.98, 2.53, 2.53, 1.31, 2.53, 1.31, 1.31, 1.31, 2.53, 2.53, 
    4.98, 1.31, 2.53, 1.31, 1.31, 2.53, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 
    1.31, 2.53, 1.31, 1.31, 2.53, 2.53, 2.53, 1.31, 2.53, 2.53, 4.98, 2.53, 
    4.98, 4.98, 6.2, 6.2, 7.42, 7.42, 12.3, 18.4, 26.95, 7.42, 6.2, 6.2, 
    7.42, 9.86, 11.08, 7.42, 8.64, 9.86, 24.51, 7.42, 6.2, 4.98, 4.98, 6.2, 
    7.42, 8.64, 8.64, 11.08, 14.74, 17.18, 17.18, 25.73, 15.96, 9.86, 7.42, 
    8.64, 2.53, 1.31, 1.31, 1.31, 1.31, 4.98, 1.31, 1.31, 1.31, 2.53, 1.31, 
    1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 
    1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 
    1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 
    1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 2.53, 1.31, 1.31, 
    1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 
    1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 2.53, 
    2.53, 1.31, 2.53, 2.53, 2.53, 4.98, 9.86, 9.86, 2.53, 2.53, 2.53, 2.53, 
    1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 2.53, 7.42, 1.31, 1.31, 1.31, 1.31, 
    1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 2.53, 4.98, 1.31, 1.31, 
    1.31, 1.31, 1.31, 1.31, 1.31, 2.53, 1.31, 2.53, 2.53, 3.75, 7.42, 22.07, 
    2.53, 2.53, 3.75, 4.98, 4.98, 7.42, 2.53, 4.98, 4.98, 7.42, 12.3, 20.84, 
    31.83, 7.42, 7.42, 7.42, 7.42, 8.64, 4.98, 1.31, 1.31, 1.31, 0.09, 1.31, 
    1.31, 1.31, 1.31, 1.31, 3.75, 7.42, 8.64, 26.95, 4.98, 4.98, 7.42, 34.27, 
    4.98, 12.3, 6.2, 7.42, 20.84, 4.98, 4.98, 15.96, 6.2, 7.42, 14.74, 36.71, 
    4.98, 1.31, 1.31, 1.31, 1.31, 2.53, 2.53, 31.83, 1.31, 1.31, 1.31, 1.31, 
    1.31, 1.31, 2.53, 4.98, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 2.53, 2.53, 
    4.98, 4.98, 9.86, 8.64, 35.49, 25.73, 12.3, 14.74, 15.96, 12.3, 12.3, 
    4.98, 3.75, 11.08, 4.98, 2.53, 2.53, 2.53, 1.31, 2.53, 1.31, 2.53, 1.31, 
    1.31, 1.31, 2.53, 1.31, 1.31, 1.31, 2.53, 4.98, 7.42, 7.42, 2.53, 2.53, 
    2.53, 1.31, 2.53, 1.31, 1.31, 4.98, 2.53, 1.31, 1.31, 1.31, 1.31, 8.64, 
    1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 
    0.09, 1.31, 1.31, 1.31, 1.31, 2.53, 1.31, 1.31, 1.31, 1.31, 1.31, 3.75, 
    3.75, 2.53, 1.31, 1.31, 2.53, 4.98, 1.31, 2.53, 1.31, 2.53, 2.53, 4.98, 
    7.42, 3.75, 2.53, 2.53, 1.31, 4.98, 2.53, 1.31, 1.31, 1.31, 1.31, 1.31, 
    2.53, 1.31, 1.31, 2.53, 2.53, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 
    1.31, 1.31, 2.53, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 2.53, 1.31, 0.09, 
    1.31, 1.31, 1.31, 2.53, 1.31, 1.31, 1.31, 2.53, 2.53, 1.31, 1.31, 3.75, 
    3.75, 1.31, 2.53, 2.53, 1.31, 1.31, 2.53, 2.53, 8.64, 6.2, 3.75, 3.75, 
    2.53, 4.98, 7.42, 1.31, 1.31, 1.31, 2.53, 4.98, 22.07, 4.98, 7.42, 31.83, 
    7.42, 12.3, 15.96, 8.64, 1.31, 2.53, 1.31, 1.31, 1.31, 2.53, 1.31, 1.31, 
    2.53, 2.53, 2.53, 2.53, 2.53, 2.53, 2.53, 7.42, 4.98, 7.42, 3.75, 4.98, 
    7.42, 18.4, 9.86, 8.64, 18.4, 6.2, 4.98, 4.98, 2.53, 4.98, 6.2, 4.98, 
    4.98, 4.98, 7.42, 7.42, 9.86, 17.18, 23.29, 11.08, 7.42, 3.75, 2.53, 
    2.53, 4.98, 1.31, 2.53, 1.31, 3.75, 1.31, 1.31, 2.53, 2.53, 1.31, 2.53, 
    6.2, 12.3, 6.2, 7.42, 36.71, 8.64, 20.84, 8.64, 12.3, 17.18, 12.3, 18.4, 
    9.86, 7.42, 8.64, 12.3, 13.52, 7.42, 18.4, 11.08, 12.3, 12.3, 12.3, 12.3, 
    12.3, 4.98, 7.42, 17.18, 11.08, 7.42, 14.74, 12.3, 1.31 ;

 TQ = 4.98, 4.98, 6.2, 6.2, 2.53, 4.98, 4.98, 4.98, 4.98, 4.98, 4.98, 4.98, 
    2.53, 3.75, 4.98, 4.98, 4.98, 6.2, 4.98, 6.2, 6.2, 20.84, 74.56, 80.66, 
    80.66, 83.1, 79.44, 79.44, 79.44, 78.22, 79.44, 77, 75.78, 75.78, 79.44, 
    79.44, 85.54, 79.44, 78.22, 85.54, 89.21, 85.54, 85.54, 86.76, 87.98, 
    89.21, 85.54, 84.32, 85.54, 90.43, 87.98, 85.54, 87.98, 90.43, 92.87, 
    94.09, 94.09, 70.89, 77, 74.56, 77, 79.44, 75.78, 75.78, 74.56, 77, 
    75.78, 85.54, 85.54, 92.87, 92.87, 87.98, 85.54, 84.32, 86.76, 89.21, 
    86.76, 85.54, 85.54, 90.43, 86.76, 90.43, 87.98, 85.54, 85.54, 90.43, 
    85.54, 83.1, 79.44, 83.1, 85.54, 73.34, 74.56, 70.89, 70.89, 70.89, 
    69.67, 70.89, 70.89, 70.89, 70.89, 69.67, 70.89, 72.12, 70.89, 73.34, 
    67.23, 70.89, 68.45, 69.67, 69.67, 66.01, 68.45, 73.34, 70.89, 68.45, 
    66.01, 70.89, 68.45, 69.67, 73.34, 70.89, 70.89, 73.34, 68.45, 70.89, 
    70.89, 73.34, 74.56, 74.56, 70.89, 70.89, 68.45, 66.01, 66.01, 66.01, 
    66.01, 67.23, 66.01, 66.01, 66.01, 68.45, 70.89, 74.56, 67.23, 79.44, 
    79.44, 84.32, 85.54, 90.43, 85.54, 85.54, 85.54, 90.43, 86.76, 80.66, 
    85.54, 85.54, 83.1, 63.57, 77, 78.22, 73.34, 74.56, 81.88, 73.34, 70.89, 
    75.78, 75.78, 79.44, 80.66, 85.54, 80.66, 83.1, 70.89, 75.78, 74.56, 
    70.89, 79.44, 79.44, 83.1, 75.78, 79.44, 79.44, 77, 70.89, 74.56, 80.66, 
    79.44, 85.54, 75.78, 69.67, 74.56, 68.45, 75.78, 75.78, 79.44, 69.67, 
    73.34, 77, 80.66, 66.01, 74.56, 74.56, 70.89, 73.34, 70.89, 74.56, 67.23, 
    70.89, 73.34, 70.89, 74.56, 86.76, 85.54, 70.89, 74.56, 74.56, 79.44, 
    83.1, 80.66, 67.23, 73.34, 77, 72.12, 77, 75.78, 77, 67.23, 63.57, 64.79, 
    64.79, 64.79, 66.01, 73.34, 74.56, 70.89, 73.34, 73.34, 73.34, 73.34, 
    70.89, 75.78, 75.78, 75.78, 83.1, 85.54, 90.43, 92.87, 92.87, 70.89, 
    73.34, 79.44, 77, 79.44, 83.1, 74.56, 79.44, 81.88, 85.54, 85.54, 94.09, 
    96.53, 95.31, 94.09, 94.09, 94.09, 85.54, 85.54, 79.44, 70.89, 63.57, 
    64.79, 77, 74.56, 77, 79.44, 83.1, 75.78, 75.78, 85.54, 77, 77, 83.1, 
    74.56, 78.22, 80.66, 74.56, 75.78, 79.44, 74.56, 74.56, 79.44, 87.98, 
    79.44, 90.43, 80.66, 94.09, 98.97, 75.78, 96.53, 79.44, 74.56, 90.43, 
    85.54, 94.09, 72.12, 77, 75.78, 74.56, 75.78, 77, 73.34, 73.34, 70.89, 
    77, 74.56, 77, 77, 74.56, 80.66, 74.56, 84.32, 83.1, 75.78, 74.56, 73.34, 
    74.56, 77, 74.56, 73.34, 74.56, 73.34, 74.56, 74.56, 72.12, 79.44, 78.22, 
    77, 78.22, 79.44, 79.44, 79.44, 79.44, 75.78, 79.44, 79.44, 77, 79.44, 
    75.78, 80.66, 80.66, 94.09, 85.54, 94.09, 92.87, 83.1, 80.66, 79.44, 
    83.1, 85.54, 94.09, 83.1, 83.1, 79.44, 74.56, 79.44, 75.78, 77, 79.44, 
    75.78, 79.44, 83.1, 79.44, 79.44, 80.66, 85.54, 90.43, 96.53, 96.53, 
    96.53, 102.63, 96.53, 105.07, 73.34, 85.54, 74.56, 91.65, 85.54, 74.56, 
    83.1, 85.54, 90.43, 79.44, 86.76, 75.78, 86.76, 77, 81.88, 79.44, 70.89, 
    73.34, 86.76, 85.54, 85.54, 85.54, 83.1, 89.21, 89.21, 86.76, 97.75, 
    90.43, 90.43, 95.31, 80.66, 85.54, 98.97, 79.44, 86.76, 90.43, 79.44, 77, 
    75.78, 83.1, 85.54, 92.87, 78.22, 79.44, 86.76, 84.32, 79.44, 75.78, 
    83.1, 77, 85.54, 73.34, 74.56, 75.78, 74.56, 86.76, 75.78, 85.54, 90.43, 
    70.89, 80.66, 86.76, 86.76, 95.31, 96.53, 94.09, 92.87, 84.32, 85.54, 
    86.76, 92.87, 85.54, 90.43, 90.43, 94.09, 102.63, 100.19, 98.97, 100.19, 
    102.63, 94.09, 101.41, 98.97, 97.75, 94.09, 98.97, 96.53, 94.09, 94.09, 
    94.09, 94.09, 101.41, 95.31, 94.09, 92.87, 98.97, 90.43, 95.31, 95.31, 
    94.09, 92.87, 86.76, 87.98, 86.76, 85.54, 85.54, 85.54, 83.1, 85.54, 
    84.32, 83.1, 85.54, 80.66, 79.44, 74.56, 80.66, 85.54, 80.66, 77, 79.44, 
    73.34, 75.78, 70.89, 77, 75.78, 79.44, 77, 79.44, 90.43, 85.54, 75.78, 
    74.56, 70.89, 75.78, 74.56, 73.34, 75.78, 75.78, 73.34, 69.67, 70.89, 
    78.22, 79.44, 86.76, 79.44, 83.1, 74.56, 85.54, 85.54, 85.54, 84.32, 
    80.66, 90.43, 85.54, 85.54, 85.54, 85.54, 85.54, 85.54, 85.54, 86.76, 
    89.21, 85.54, 86.76, 87.98, 85.54, 85.54, 79.44, 79.44, 81.88, 80.66, 
    83.1, 80.66, 81.88, 80.66, 84.32, 83.1, 79.44, 79.44, 85.54, 79.44, 
    79.44, 78.22, 80.66, 81.88, 80.66, 79.44, 79.44, 80.66, 79.44, 77, 80.66, 
    79.44, 79.44, 79.44, 81.88, 85.54, 79.44, 84.32, 83.1, 83.1, 79.44, 
    80.66, 84.32, 80.66, 84.32, 79.44, 79.44, 79.44, 83.1, 85.54, 85.54, 
    90.43, 92.87, 87.98, 86.76, 86.76, 84.32, 90.43, 85.54, 85.54, 84.32, 
    83.1, 83.1, 85.54, 85.54, 94.09, 92.87, 94.09, 85.54, 83.1, 86.76, 74.56, 
    81.88, 79.44, 80.66, 98.97, 86.76, 83.1, 90.43, 87.98, 85.54, 98.97, 
    103.85, 94.09, 85.54, 85.54, 85.54, 79.44, 78.22, 75.78, 75.78, 79.44, 
    85.54, 86.76, 89.21, 98.97, 83.1, 81.88, 80.66, 85.54, 79.44, 90.43, 
    90.43, 92.87, 95.31, 90.43, 90.43, 85.54, 94.09, 90.43, 92.87, 74.56, 
    85.54, 97.75, 98.97, 85.54, 94.09, 90.43, 79.44, 92.87, 96.53, 90.43, 
    83.1, 81.88, 78.22, 80.66, 90.43, 90.43, 94.09, 83.1, 73.34, 78.22, 77, 
    79.44, 80.66, 85.54, 94.09, 97.75, 98.97, 92.87, 96.53, 89.21, 90.43, 
    81.88, 85.54, 86.76, 94.09, 78.22, 81.88, 85.54, 79.44, 89.21, 86.76, 
    83.1, 85.54, 85.54, 72.12, 85.54, 86.76, 69.67, 77, 83.1, 85.54, 92.87, 
    80.66, 80.66, 85.54, 64.79, 85.54, 98.97, 86.76, 85.54, 80.66, 83.1, 
    89.21, 78.22, 79.44, 79.44, 85.54, 90.43, 92.87, 85.54, 83.1, 81.88, 
    84.32, 80.66, 75.78, 74.56, 61.13, 64.79, 74.56, 84.32, 78.22, 79.44, 
    85.54, 85.54, 85.54, 70.89, 74.56, 77, 77, 74.56, 79.44, 75.78, 78.22, 
    80.66, 79.44, 80.66, 77, 78.22, 80.66, 79.44, 83.1, 80.66, 79.44, 77, 
    75.78, 79.44, 79.44, 79.44, 83.1, 85.54, 90.43, 79.44, 83.1, 74.56, 77, 
    79.44, 86.76, 79.44, 75.78, 75.78, 75.78, 77, 77, 75.78, 75.78, 74.56, 
    74.56, 75.78, 74.56, 77, 77, 77, 79.44, 73.34, 77, 87.98, 79.44, 81.88, 
    85.54, 80.66, 79.44, 90.43, 92.87, 74.56, 77, 79.44, 78.22, 85.54, 73.34, 
    79.44, 80.66, 79.44, 80.66, 84.32, 89.21, 70.89, 79.44, 80.66, 80.66, 
    79.44, 83.1, 77, 79.44, 79.44, 83.1, 79.44, 83.1, 79.44, 79.44, 79.44, 
    79.44, 106.3, 89.21, 77, 75.78, 83.1, 74.56, 79.44, 73.34, 74.56, 74.56, 
    77, 78.22, 74.56, 75.78, 77, 77, 75.78, 78.22, 73.34, 70.89, 74.56, 
    74.56, 75.78, 70.89, 70.89, 79.44, 77, 81.88, 90.43, 74.56, 77, 90.43, 
    79.44, 79.44, 79.44, 79.44, 80.66, 77, 85.54, 85.54, 85.54, 77, 86.76, 
    83.1, 86.76, 92.87, 83.1, 74.56, 85.54, 90.43, 91.65, 90.43, 85.54, 
    84.32, 89.21, 69.67, 86.76, 85.54, 78.22, 79.44, 73.34, 74.56, 75.78, 
    74.56, 70.89, 74.56, 75.78, 77, 89.21, 85.54, 81.88, 79.44, 79.44, 83.1, 
    83.1, 83.1, 77, 75.78, 83.1, 77, 86.76, 74.56, 83.1, 78.22, 77, 77, 77, 
    83.1, 79.44, 75.78, 78.22, 86.76, 80.66, 79.44, 84.32, 83.1, 83.1, 80.66, 
    77, 73.34, 77, 75.78, 74.56, 75.78, 75.78, 79.44, 74.56, 75.78, 70.89, 
    77, 94.09, 79.44, 84.32, 87.98, 92.87, 96.53, 80.66, 75.78, 77, 67.23, 
    74.56, 75.78, 74.56, 70.89, 70.89, 75.78, 74.56, 77, 79.44, 83.1, 73.34, 
    79.44, 77, 85.54, 86.76, 92.87, 85.54, 77, 84.32, 79.44, 75.78, 83.1, 77, 
    74.56, 86.76, 85.54, 85.54, 64.79 ;

 SP = 1.31, 2.53, 1.31, 0, 4.98, 1.31, 0.09, 1.31, 6.2, 0, 4.98, 1.31, 2.53, 
    2.53, 1.31, 1.31, 2.53, 1.31, 1.31, 1.31, 2.53, 2.53, 1.31, 2.53, 0.09, 
    0, 1.31, 4.98, 2.53, 2.53, 1.31, 1.31, 4.98, 0, 1.31, 2.53, 4.98, 4.98, 
    0, 0.09, 2.53, 1.31, 2.53, 1.31, 1.31, 1.31, 0, 1.31, 1.31, 4.98, 1.31, 
    1.31, 1.31, 0, 1.31, 1.31, 0, 4.98, 4.98, 1.31, 1.31, 1.31, 2.53, 2.53, 
    2.53, 4.98, 1.31, 1.31, 2.53, 0, 1.31, 2.53, 1.31, 1.31, 1.31, 1.31, 
    1.31, 2.53, 0, 2.53, 0, 4.98, 1.31, 2.53, 4.98, 2.53, 1.31, 1.31, 2.53, 
    0, 1.31, 1.31, 6.2, 4.98, 2.53, 3.75, 1.31, 0, 2.53, 0, 1.31, 0, 1.31, 
    1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 6.2, 1.31, 0, 2.53, 4.98, 1.31, 
    1.31, 0, 1.31, 1.31, 2.53, 1.31, 2.53, 2.53, 1.31, 2.53, 1.31, 1.31, 0, 
    2.53, 1.31, 4.98, 1.31, 2.53, 2.53, 2.53, 2.53, 0, 1.31, 2.53, 1.31, 
    1.31, 2.53, 4.98, 1.31, 1.31, 0, 2.53, 1.31, 1.31, 1.31, 2.53, 1.31, 
    4.98, 1.31, 1.31, 2.53, 0, 2.53, 6.2, 6.2, 2.53, 2.53, 6.2, 1.31, 2.53, 
    2.53, 6.2, 1.31, 4.98, 1.31, 4.98, 3.75, 2.53, 1.31, 1.31, 1.31, 6.2, 
    2.53, 1.31, 2.53, 4.98, 2.53, 2.53, 1.31, 1.31, 2.53, 4.98, 4.98, 0.09, 
    2.53, 3.75, 1.31, 4.98, 1.31, 2.53, 0, 2.53, 4.98, 0, 1.31, 2.53, 3.75, 
    1.31, 4.98, 2.53, 2.53, 1.31, 6.2, 4.98, 1.31, 4.98, 1.31, 1.31, 1.31, 
    4.98, 1.31, 0, 2.53, 4.98, 1.31, 1.31, 1.31, 2.53, 0, 2.53, 0, 6.2, 1.31, 
    2.53, 1.31, 6.2, 7.42, 0, 2.53, 1.31, 4.98, 1.31, 1.31, 2.53, 2.53, 6.2, 
    0, 1.31, 1.31, 4.98, 4.98, 4.98, 0, 1.31, 6.2, 2.53, 3.75, 1.31, 4.98, 
    1.31, 4.98, 2.53, 1.31, 1.31, 4.98, 2.53, 2.53, 0, 1.31, 2.53, 0, 2.53, 
    2.53, 4.98, 4.98, 3.75, 2.53, 1.31, 4.98, 1.31, 4.98, 2.53, 1.31, 1.31, 
    2.53, 2.53, 4.98, 2.53, 2.53, 1.31, 1.31, 0, 2.53, 2.53, 0, 1.31, 2.53, 
    4.98, 1.31, 1.31, 3.75, 1.31, 4.98, 2.53, 4.98, 1.31, 2.53, 1.31, 0, 
    2.53, 3.75, 4.98, 2.53, 2.53, 0.09, 6.2, 1.31, 2.53, 4.98, 1.31, 2.53, 
    4.98, 1.31, 1.31, 4.98, 1.31, 2.53, 1.31, 1.31, 2.53, 1.31, 1.31, 1.31, 
    2.53, 1.31, 3.75, 4.98, 6.2, 0, 1.31, 1.31, 2.53, 4.98, 4.98, 1.31, 0, 
    4.98, 2.53, 4.98, 1.31, 4.98, 1.31, 1.31, 6.2, 3.75, 2.53, 6.2, 6.2, 
    1.31, 1.31, 1.31, 3.75, 1.31, 1.31, 2.53, 1.31, 0, 6.2, 2.53, 4.98, 2.53, 
    1.31, 0, 0, 1.31, 2.53, 4.98, 6.2, 1.31, 7.42, 1.31, 1.31, 2.53, 2.53, 
    1.31, 1.31, 2.53, 1.31, 1.31, 1.31, 4.98, 2.53, 4.98, 6.2, 1.31, 1.31, 
    1.31, 6.2, 2.53, 4.98, 4.98, 6.2, 0, 2.53, 0, 2.53, 6.2, 4.98, 1.31, 
    1.31, 4.98, 2.53, 3.75, 6.2, 0, 4.98, 1.31, 1.31, 2.53, 1.31, 1.31, 4.98, 
    4.98, 4.98, 1.31, 6.2, 2.53, 1.31, 1.31, 4.98, 2.53, 0, 1.31, 2.53, 1.31, 
    1.31, 2.53, 7.42, 3.75, 6.2, 2.53, 2.53, 1.31, 1.31, 2.53, 4.98, 2.53, 
    2.53, 0.09, 2.53, 0.09, 3.75, 3.75, 4.98, 1.31, 2.53, 1.31, 2.53, 1.31, 
    6.2, 1.31, 1.31, 2.53, 2.53, 2.53, 6.2, 0, 1.31, 1.31, 4.98, 2.53, 6.2, 
    4.98, 1.31, 1.31, 1.31, 2.53, 4.98, 1.31, 1.31, 0, 4.98, 2.53, 3.75, 
    1.31, 1.31, 2.53, 4.98, 4.98, 1.31, 1.31, 1.31, 6.2, 2.53, 4.98, 0, 2.53, 
    0, 6.2, 1.31, 1.31, 2.53, 1.31, 2.53, 1.31, 1.31, 3.75, 0, 3.75, 1.31, 
    2.53, 2.53, 1.31, 1.31, 0, 4.98, 2.53, 1.31, 2.53, 1.31, 6.2, 1.31, 1.31, 
    2.53, 4.98, 2.53, 2.53, 4.98, 1.31, 6.2, 2.53, 7.42, 4.98, 1.31, 2.53, 
    2.53, 1.31, 1.31, 4.98, 0.09, 1.31, 1.31, 0.09, 2.53, 4.98, 0, 1.31, 
    1.31, 0, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 1.31, 0, 1.31, 
    1.31, 1.31, 3.75, 1.31, 1.31, 4.98, 0, 1.31, 1.31, 2.53, 2.53, 1.31, 
    1.31, 1.31, 2.53, 4.98, 4.98, 0.09, 0, 1.31, 1.31, 1.31, 1.31, 1.31, 
    1.31, 1.31, 3.75, 0, 1.31, 2.53, 1.31, 4.98, 1.31, 2.53, 0, 1.31, 1.31, 
    2.53, 2.53, 6.2, 3.75, 2.53, 0, 2.53, 4.98, 4.98, 2.53, 1.31, 2.53, 2.53, 
    2.53, 2.53, 1.31, 2.53, 7.42, 3.75, 3.75, 6.2, 1.31, 4.98, 3.75, 2.53, 
    4.98, 1.31, 1.31, 0, 4.98, 1.31, 3.75, 3.75, 2.53, 4.98, 1.31, 4.98, 
    4.98, 1.31, 2.53, 1.31, 2.53, 1.31, 2.53, 2.53, 1.31, 2.53, 1.31, 2.53, 
    1.31, 2.53, 2.53, 1.31, 1.31, 2.53, 1.31, 2.53, 2.53, 1.31, 2.53, 2.53, 
    4.98, 1.31, 1.31, 2.53, 2.53, 2.53, 4.98, 1.31, 0, 2.53, 2.53, 1.31, 
    2.53, 1.31, 2.53, 1.31, 3.75, 4.98, 3.75, 4.98, 0, 2.53, 1.31, 1.31, 
    1.31, 3.75, 1.31, 1.31, 2.53, 2.53, 2.53, 3.75, 1.31, 1.31, 1.31, 1.31, 
    4.98, 2.53, 4.98, 1.31, 2.53, 2.53, 1.31, 2.53, 1.31, 1.31, 1.31, 1.31, 
    4.98, 2.53, 4.98, 4.98, 1.31, 2.53, 0, 0.09, 1.31, 0, 0, 1.31, 3.75, 0, 
    0, 0, 2.53, 1.31, 4.98, 4.98, 2.53, 2.53, 1.31, 2.53, 2.53, 4.98, 4.98, 
    4.98, 4.98, 1.31, 2.53, 2.53, 1.31, 2.53, 0, 2.53, 1.31, 0, 1.31, 2.53, 
    1.31, 4.98, 2.53, 1.31, 1.31, 1.31, 1.31, 0.09, 1.31, 2.53, 4.98, 1.31, 
    4.98, 4.98, 0, 1.31, 6.2, 4.98, 4.98, 4.98, 1.31, 1.31, 1.31, 1.31, 4.98, 
    0, 2.53, 2.53, 2.53, 1.31, 4.98, 1.31, 2.53, 2.53, 2.53, 1.31, 2.53, 
    4.98, 1.31, 2.53, 2.53, 4.98, 2.53, 4.98, 1.31, 2.53, 1.31, 2.53, 1.31, 
    1.31, 1.31, 1.31, 2.53, 7.42, 2.53, 2.53, 0.09, 2.53, 2.53, 7.42, 4.98, 
    2.53, 1.31, 0, 2.53, 2.53, 1.31, 1.31, 1.31, 1.31, 1.31, 6.2, 3.75, 1.31, 
    1.31, 2.53, 2.53, 1.31, 0, 1.31, 1.31, 2.53, 4.98, 1.31, 4.98, 1.31, 
    2.53, 2.53, 7.42, 0.09, 6.2, 0, 2.53, 1.31, 2.53, 2.53, 4.98, 4.98, 2.53, 
    0, 0, 0, 1.31, 2.53, 1.31, 1.31, 0, 0.09, 2.53, 1.31, 1.31, 2.53, 2.53, 
    2.53, 2.53, 4.98, 2.53, 2.53, 2.53, 1.31, 2.53, 1.31, 1.31, 4.98, 2.53, 
    4.98, 1.31, 2.53, 3.75, 1.31, 4.98, 1.31, 2.53, 3.75, 1.31, 2.53, 2.53, 
    2.53, 0, 1.31, 1.31, 4.98, 4.98, 7.42, 4.98, 1.31, 0, 1.31, 3.75, 2.53, 
    2.53, 3.75, 2.53, 1.31, 1.31, 2.53, 1.31, 6.2, 4.98, 1.31, 1.31, 4.98, 
    4.98, 3.75, 2.53, 6.2, 2.53, 1.31, 1.31, 4.98, 2.53, 2.53, 3.75, 6.2, 
    2.53, 1.31, 3.75, 1.31, 2.53, 6.2, 4.98, 2.53, 2.53, 2.53, 1.31, 2.53, 
    1.31, 1.31, 1.31, 2.53, 2.53, 1.31, 0, 1.31, 2.53, 2.53, 6.2, 0, 0, 1.31, 
    6.2, 2.53, 1.31, 2.53, 1.31, 1.31, 2.53, 6.2, 1.31, 0.09, 1.31, 2.53, 
    2.53, 1.31, 2.53, 3.75, 1.31, 3.75, 1.31, 2.53, 4.98, 1.31, 2.53, 1.31, 
    2.53, 1.31, 2.53, 1.31, 2.53, 4.98, 0, 4.98, 4.98, 7.42 ;
}
